module rvclkhdr(
  output  io_l1clk,
  input   io_clk,
  input   io_en,
  input   io_scan_mode
);
  wire  clkhdr_Q; // @[el2_lib.scala 474:26]
  wire  clkhdr_CK; // @[el2_lib.scala 474:26]
  wire  clkhdr_EN; // @[el2_lib.scala 474:26]
  wire  clkhdr_SE; // @[el2_lib.scala 474:26]
  gated_latch clkhdr ( // @[el2_lib.scala 474:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign io_l1clk = clkhdr_Q; // @[el2_lib.scala 475:14]
  assign clkhdr_CK = io_clk; // @[el2_lib.scala 476:18]
  assign clkhdr_EN = io_en; // @[el2_lib.scala 477:18]
  assign clkhdr_SE = io_scan_mode; // @[el2_lib.scala 478:18]
endmodule
module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [63:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [63:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_scan_mode; // @[el2_lib.scala 483:22]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 186:53]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 322:61]
  wire  _T_319 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 323:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_319; // @[el2_ifu_mem_ctl.scala 323:42]
  wire  _T = io_ifc_fetch_req_bf_raw | ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 187:53]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 254:30]
  wire  _T_1 = _T | miss_pending; // @[el2_ifu_mem_ctl.scala 187:71]
  wire  _T_2 = _T_1 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 187:86]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 552:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_319; // @[el2_ifu_mem_ctl.scala 554:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 188:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 309:63]
  wire [4:0] _GEN_437 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 670:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_437 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 670:53]
  wire [1:0] _GEN_438 = {{1'd0}, _T_319}; // @[el2_ifu_mem_ctl.scala 673:91]
  wire [1:0] _T_3080 = ic_fetch_val_shift_right[3:2] & _GEN_438; // @[el2_ifu_mem_ctl.scala 673:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 324:60]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 276:46]
  wire [1:0] _GEN_439 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 673:113]
  wire [1:0] _T_3081 = _T_3080 & _GEN_439; // @[el2_ifu_mem_ctl.scala 673:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 659:59]
  wire [1:0] _GEN_440 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 673:130]
  wire [1:0] _T_3082 = _T_3081 | _GEN_440; // @[el2_ifu_mem_ctl.scala 673:130]
  wire  _T_3083 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 673:154]
  wire [1:0] _GEN_441 = {{1'd0}, _T_3083}; // @[el2_ifu_mem_ctl.scala 673:152]
  wire [1:0] _T_3084 = _T_3082 & _GEN_441; // @[el2_ifu_mem_ctl.scala 673:152]
  wire [1:0] _T_3073 = ic_fetch_val_shift_right[1:0] & _GEN_438; // @[el2_ifu_mem_ctl.scala 673:91]
  wire [1:0] _T_3074 = _T_3073 & _GEN_439; // @[el2_ifu_mem_ctl.scala 673:113]
  wire [1:0] _T_3075 = _T_3074 | _GEN_440; // @[el2_ifu_mem_ctl.scala 673:130]
  wire [1:0] _T_3077 = _T_3075 & _GEN_441; // @[el2_ifu_mem_ctl.scala 673:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3084,_T_3077}; // @[Cat.scala 29:58]
  wire  _T_3184 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 333:30]
  wire  _T_3185 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 333:44]
  wire  _T_3186 = _T_3184 ^ _T_3185; // @[el2_lib.scala 333:35]
  wire [5:0] _T_3194 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 333:76]
  wire  _T_3195 = ^_T_3194; // @[el2_lib.scala 333:83]
  wire  _T_3196 = io_iccm_rd_data_ecc[37] ^ _T_3195; // @[el2_lib.scala 333:71]
  wire [6:0] _T_3203 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 333:103]
  wire [14:0] _T_3211 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3203}; // @[el2_lib.scala 333:103]
  wire  _T_3212 = ^_T_3211; // @[el2_lib.scala 333:110]
  wire  _T_3213 = io_iccm_rd_data_ecc[36] ^ _T_3212; // @[el2_lib.scala 333:98]
  wire [6:0] _T_3220 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 333:130]
  wire [14:0] _T_3228 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3220}; // @[el2_lib.scala 333:130]
  wire  _T_3229 = ^_T_3228; // @[el2_lib.scala 333:137]
  wire  _T_3230 = io_iccm_rd_data_ecc[35] ^ _T_3229; // @[el2_lib.scala 333:125]
  wire [8:0] _T_3239 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 333:157]
  wire [17:0] _T_3248 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3239}; // @[el2_lib.scala 333:157]
  wire  _T_3249 = ^_T_3248; // @[el2_lib.scala 333:164]
  wire  _T_3250 = io_iccm_rd_data_ecc[34] ^ _T_3249; // @[el2_lib.scala 333:152]
  wire [8:0] _T_3259 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 333:184]
  wire [17:0] _T_3268 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3259}; // @[el2_lib.scala 333:184]
  wire  _T_3269 = ^_T_3268; // @[el2_lib.scala 333:191]
  wire  _T_3270 = io_iccm_rd_data_ecc[33] ^ _T_3269; // @[el2_lib.scala 333:179]
  wire [8:0] _T_3279 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 333:211]
  wire [17:0] _T_3288 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3279}; // @[el2_lib.scala 333:211]
  wire  _T_3289 = ^_T_3288; // @[el2_lib.scala 333:218]
  wire  _T_3290 = io_iccm_rd_data_ecc[32] ^ _T_3289; // @[el2_lib.scala 333:206]
  wire [6:0] _T_3296 = {_T_3186,_T_3196,_T_3213,_T_3230,_T_3250,_T_3270,_T_3290}; // @[Cat.scala 29:58]
  wire  _T_3297 = _T_3296 != 7'h0; // @[el2_lib.scala 334:44]
  wire  _T_3298 = iccm_ecc_word_enable[0] & _T_3297; // @[el2_lib.scala 334:32]
  wire  _T_3300 = _T_3298 & _T_3296[6]; // @[el2_lib.scala 334:53]
  wire  _T_3569 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 333:30]
  wire  _T_3570 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 333:44]
  wire  _T_3571 = _T_3569 ^ _T_3570; // @[el2_lib.scala 333:35]
  wire [5:0] _T_3579 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 333:76]
  wire  _T_3580 = ^_T_3579; // @[el2_lib.scala 333:83]
  wire  _T_3581 = io_iccm_rd_data_ecc[76] ^ _T_3580; // @[el2_lib.scala 333:71]
  wire [6:0] _T_3588 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 333:103]
  wire [14:0] _T_3596 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3588}; // @[el2_lib.scala 333:103]
  wire  _T_3597 = ^_T_3596; // @[el2_lib.scala 333:110]
  wire  _T_3598 = io_iccm_rd_data_ecc[75] ^ _T_3597; // @[el2_lib.scala 333:98]
  wire [6:0] _T_3605 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 333:130]
  wire [14:0] _T_3613 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3605}; // @[el2_lib.scala 333:130]
  wire  _T_3614 = ^_T_3613; // @[el2_lib.scala 333:137]
  wire  _T_3615 = io_iccm_rd_data_ecc[74] ^ _T_3614; // @[el2_lib.scala 333:125]
  wire [8:0] _T_3624 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 333:157]
  wire [17:0] _T_3633 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3624}; // @[el2_lib.scala 333:157]
  wire  _T_3634 = ^_T_3633; // @[el2_lib.scala 333:164]
  wire  _T_3635 = io_iccm_rd_data_ecc[73] ^ _T_3634; // @[el2_lib.scala 333:152]
  wire [8:0] _T_3644 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 333:184]
  wire [17:0] _T_3653 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3644}; // @[el2_lib.scala 333:184]
  wire  _T_3654 = ^_T_3653; // @[el2_lib.scala 333:191]
  wire  _T_3655 = io_iccm_rd_data_ecc[72] ^ _T_3654; // @[el2_lib.scala 333:179]
  wire [8:0] _T_3664 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 333:211]
  wire [17:0] _T_3673 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3664}; // @[el2_lib.scala 333:211]
  wire  _T_3674 = ^_T_3673; // @[el2_lib.scala 333:218]
  wire  _T_3675 = io_iccm_rd_data_ecc[71] ^ _T_3674; // @[el2_lib.scala 333:206]
  wire [6:0] _T_3681 = {_T_3571,_T_3581,_T_3598,_T_3615,_T_3635,_T_3655,_T_3675}; // @[Cat.scala 29:58]
  wire  _T_3682 = _T_3681 != 7'h0; // @[el2_lib.scala 334:44]
  wire  _T_3683 = iccm_ecc_word_enable[1] & _T_3682; // @[el2_lib.scala 334:32]
  wire  _T_3685 = _T_3683 & _T_3681[6]; // @[el2_lib.scala 334:53]
  wire [1:0] iccm_single_ecc_error = {_T_3300,_T_3685}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 191:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 636:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 192:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 193:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 479:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 193:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 193:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 193:72]
  wire  _T_2477 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2482 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2502 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 529:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 392:42]
  wire  _T_2504 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 529:79]
  wire  _T_2505 = _T_2502 | _T_2504; // @[el2_ifu_mem_ctl.scala 529:56]
  wire  _T_2506 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 529:122]
  wire  _T_2507 = ~_T_2506; // @[el2_ifu_mem_ctl.scala 529:101]
  wire  _T_2508 = _T_2505 & _T_2507; // @[el2_ifu_mem_ctl.scala 529:99]
  wire  _T_2509 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2523 = io_ifu_fetch_val[0] & _T_319; // @[el2_ifu_mem_ctl.scala 536:45]
  wire  _T_2524 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 536:69]
  wire  _T_2525 = _T_2523 & _T_2524; // @[el2_ifu_mem_ctl.scala 536:67]
  wire  _T_2526 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_2509 ? _T_2525 : _T_2526; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2482 ? _T_2508 : _GEN_38; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2477 ? 1'h0 : _GEN_42; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 193:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 195:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 195:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 284:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 284:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 705:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 284:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 275:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 275:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 326:71]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 275:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 275:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 284:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 284:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 284:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 284:114]
  reg  ifu_bus_rvalid_unq_ff; // @[el2_ifu_mem_ctl.scala 579:56]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 551:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 593:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 620:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 311:62]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 601:56]
  wire  _T_2623 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 618:69]
  wire  _T_2624 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 618:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2623 : _T_2624; // @[el2_ifu_mem_ctl.scala 618:28]
  wire  _T_2575 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 597:68]
  wire  _T_2576 = ic_act_miss_f | _T_2575; // @[el2_ifu_mem_ctl.scala 597:48]
  wire  bus_reset_data_beat_cnt = _T_2576 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 597:91]
  wire  _T_2572 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 596:50]
  wire  _T_2573 = bus_ifu_wr_en_ff & _T_2572; // @[el2_ifu_mem_ctl.scala 596:48]
  wire  _T_2574 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 596:72]
  wire  bus_inc_data_beat_cnt = _T_2573 & _T_2574; // @[el2_ifu_mem_ctl.scala 596:70]
  wire [2:0] _T_2580 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 600:115]
  wire [2:0] _T_2582 = bus_inc_data_beat_cnt ? _T_2580 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2577 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 598:32]
  wire  _T_2578 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 598:57]
  wire  bus_hold_data_beat_cnt = _T_2577 & _T_2578; // @[el2_ifu_mem_ctl.scala 598:55]
  wire [2:0] _T_2583 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2582 | _T_2583; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 195:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 195:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 196:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 195:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 196:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_319; // @[el2_ifu_mem_ctl.scala 202:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 202:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 429:45]
  wire  _T_2106 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 450:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 406:60]
  wire  _T_2137 = _T_2106 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2110 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 450:127]
  wire  _T_2138 = _T_2110 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2145 = _T_2137 | _T_2138; // @[Mux.scala 27:72]
  wire  _T_2114 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 450:127]
  wire  _T_2139 = _T_2114 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2146 = _T_2145 | _T_2139; // @[Mux.scala 27:72]
  wire  _T_2118 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 450:127]
  wire  _T_2140 = _T_2118 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2147 = _T_2146 | _T_2140; // @[Mux.scala 27:72]
  wire  _T_2122 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 450:127]
  wire  _T_2141 = _T_2122 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2148 = _T_2147 | _T_2141; // @[Mux.scala 27:72]
  wire  _T_2126 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 450:127]
  wire  _T_2142 = _T_2126 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2149 = _T_2148 | _T_2142; // @[Mux.scala 27:72]
  wire  _T_2130 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 450:127]
  wire  _T_2143 = _T_2130 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2150 = _T_2149 | _T_2143; // @[Mux.scala 27:72]
  wire  _T_2134 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 450:127]
  wire  _T_2144 = _T_2134 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2150 | _T_2144; // @[Mux.scala 27:72]
  wire  _T_2192 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 452:69]
  wire  _T_2193 = ic_miss_buff_data_valid_bypass_index & _T_2192; // @[el2_ifu_mem_ctl.scala 452:67]
  wire  _T_2195 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 452:91]
  wire  _T_2196 = _T_2193 & _T_2195; // @[el2_ifu_mem_ctl.scala 452:89]
  wire  _T_2201 = _T_2193 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 453:65]
  wire  _T_2202 = _T_2196 | _T_2201; // @[el2_ifu_mem_ctl.scala 452:112]
  wire  _T_2204 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 454:43]
  wire  _T_2207 = _T_2204 & _T_2195; // @[el2_ifu_mem_ctl.scala 454:65]
  wire  _T_2208 = _T_2202 | _T_2207; // @[el2_ifu_mem_ctl.scala 453:88]
  wire  _T_2212 = _T_2204 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 455:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 432:75]
  wire  _T_2152 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 451:110]
  wire  _T_2176 = _T_2152 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2155 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 451:110]
  wire  _T_2177 = _T_2155 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2184 = _T_2176 | _T_2177; // @[Mux.scala 27:72]
  wire  _T_2158 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 451:110]
  wire  _T_2178 = _T_2158 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2185 = _T_2184 | _T_2178; // @[Mux.scala 27:72]
  wire  _T_2161 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 451:110]
  wire  _T_2179 = _T_2161 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2186 = _T_2185 | _T_2179; // @[Mux.scala 27:72]
  wire  _T_2164 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 451:110]
  wire  _T_2180 = _T_2164 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2187 = _T_2186 | _T_2180; // @[Mux.scala 27:72]
  wire  _T_2167 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 451:110]
  wire  _T_2181 = _T_2167 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2188 = _T_2187 | _T_2181; // @[Mux.scala 27:72]
  wire  _T_2170 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 451:110]
  wire  _T_2182 = _T_2170 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2189 = _T_2188 | _T_2182; // @[Mux.scala 27:72]
  wire  _T_2173 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 451:110]
  wire  _T_2183 = _T_2173 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2189 | _T_2183; // @[Mux.scala 27:72]
  wire  _T_2213 = _T_2212 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 455:87]
  wire  _T_2214 = _T_2208 | _T_2213; // @[el2_ifu_mem_ctl.scala 454:88]
  wire  _T_2218 = ic_miss_buff_data_valid_bypass_index & _T_2134; // @[el2_ifu_mem_ctl.scala 456:43]
  wire  miss_buff_hit_unq_f = _T_2214 | _T_2218; // @[el2_ifu_mem_ctl.scala 455:131]
  wire  _T_2234 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 461:55]
  wire  _T_2235 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 461:87]
  wire  _T_2236 = _T_2234 | _T_2235; // @[el2_ifu_mem_ctl.scala 461:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2236; // @[el2_ifu_mem_ctl.scala 461:41]
  wire  _T_2219 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 458:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 312:49]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[el2_ifu_mem_ctl.scala 449:51]
  wire  _T_2220 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 458:68]
  wire  _T_2221 = miss_buff_hit_unq_f & _T_2220; // @[el2_ifu_mem_ctl.scala 458:66]
  wire  stream_hit_f = _T_2219 & _T_2221; // @[el2_ifu_mem_ctl.scala 458:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 279:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 279:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 279:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 603:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 630:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 206:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 206:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 206:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 206:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 207:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 207:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 207:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 208:16]
  wire  _T_44 = _T_42 & _T_319; // @[el2_ifu_mem_ctl.scala 208:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 208:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 208:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 209:49]
  wire  _T_54 = ic_byp_hit_f & _T_319; // @[el2_ifu_mem_ctl.scala 210:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 210:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 210:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 198:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 210:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 210:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 210:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_319; // @[el2_ifu_mem_ctl.scala 211:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 211:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 211:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 211:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 212:102]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 213:46]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 213:70]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 213:24]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 212:22]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 211:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 210:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 209:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 208:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 207:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 206:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2231 = byp_fetch_index[4:1] == 4'hf; // @[el2_ifu_mem_ctl.scala 460:60]
  wire  _T_2232 = _T_2231 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 460:94]
  wire  stream_eol_f = _T_2232 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 460:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 221:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 221:87]
  wire  _T_113 = _T_111 & _T_2574; // @[el2_ifu_mem_ctl.scala 221:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 221:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 225:48]
  wire  _T_126 = _T_124 & _T_2574; // @[el2_ifu_mem_ctl.scala 225:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 225:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 285:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 285:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 285:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 285:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 285:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 286:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 285:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 286:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 340:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 286:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 286:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 286:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 229:50]
  wire  _T_137 = _T_135 & _T_2574; // @[el2_ifu_mem_ctl.scala 229:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 287:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 288:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 288:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 287:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 230:35]
  wire  _T_143 = _T_141 & _T_2574; // @[el2_ifu_mem_ctl.scala 230:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 230:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 229:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 235:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 234:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 234:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 239:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 239:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 196:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 196:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 196:26]
  wire  _T_30 = ic_act_miss_f & _T_2574; // @[el2_ifu_mem_ctl.scala 203:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 214:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 214:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 214:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 214:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 214:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 214:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 218:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 218:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 218:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 222:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 222:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 226:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 226:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 231:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 231:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 231:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 236:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 236:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 255:95]
  wire  _T_175 = _T_2234 & _T_174; // @[el2_ifu_mem_ctl.scala 255:93]
  wire  crit_wd_byp_ok_ff = _T_2235 | _T_175; // @[el2_ifu_mem_ctl.scala 255:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 256:36]
  wire  _T_180 = _T_2234 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 256:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 256:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 256:70]
  wire  _T_184 = _T_2234 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 257:39]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 257:5]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 256:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 257:59]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 258:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 258:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 257:75]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 260:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 260:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:64]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[el2_ifu_mem_ctl.scala 737:12]
  wire  _T_4620 = ifu_ic_rw_int_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire  _T_4748 = _T_4620 & way_status_out_0; // @[Mux.scala 27:72]
  wire  _T_4621 = ifu_ic_rw_int_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire  _T_4749 = _T_4621 & way_status_out_1; // @[Mux.scala 27:72]
  wire  _T_4876 = _T_4748 | _T_4749; // @[Mux.scala 27:72]
  wire  _T_4622 = ifu_ic_rw_int_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire  _T_4750 = _T_4622 & way_status_out_2; // @[Mux.scala 27:72]
  wire  _T_4877 = _T_4876 | _T_4750; // @[Mux.scala 27:72]
  wire  _T_4623 = ifu_ic_rw_int_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire  _T_4751 = _T_4623 & way_status_out_3; // @[Mux.scala 27:72]
  wire  _T_4878 = _T_4877 | _T_4751; // @[Mux.scala 27:72]
  wire  _T_4624 = ifu_ic_rw_int_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire  _T_4752 = _T_4624 & way_status_out_4; // @[Mux.scala 27:72]
  wire  _T_4879 = _T_4878 | _T_4752; // @[Mux.scala 27:72]
  wire  _T_4625 = ifu_ic_rw_int_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire  _T_4753 = _T_4625 & way_status_out_5; // @[Mux.scala 27:72]
  wire  _T_4880 = _T_4879 | _T_4753; // @[Mux.scala 27:72]
  wire  _T_4626 = ifu_ic_rw_int_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire  _T_4754 = _T_4626 & way_status_out_6; // @[Mux.scala 27:72]
  wire  _T_4881 = _T_4880 | _T_4754; // @[Mux.scala 27:72]
  wire  _T_4627 = ifu_ic_rw_int_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire  _T_4755 = _T_4627 & way_status_out_7; // @[Mux.scala 27:72]
  wire  _T_4882 = _T_4881 | _T_4755; // @[Mux.scala 27:72]
  wire  _T_4628 = ifu_ic_rw_int_addr_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire  _T_4756 = _T_4628 & way_status_out_8; // @[Mux.scala 27:72]
  wire  _T_4883 = _T_4882 | _T_4756; // @[Mux.scala 27:72]
  wire  _T_4629 = ifu_ic_rw_int_addr_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire  _T_4757 = _T_4629 & way_status_out_9; // @[Mux.scala 27:72]
  wire  _T_4884 = _T_4883 | _T_4757; // @[Mux.scala 27:72]
  wire  _T_4630 = ifu_ic_rw_int_addr_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire  _T_4758 = _T_4630 & way_status_out_10; // @[Mux.scala 27:72]
  wire  _T_4885 = _T_4884 | _T_4758; // @[Mux.scala 27:72]
  wire  _T_4631 = ifu_ic_rw_int_addr_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire  _T_4759 = _T_4631 & way_status_out_11; // @[Mux.scala 27:72]
  wire  _T_4886 = _T_4885 | _T_4759; // @[Mux.scala 27:72]
  wire  _T_4632 = ifu_ic_rw_int_addr_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire  _T_4760 = _T_4632 & way_status_out_12; // @[Mux.scala 27:72]
  wire  _T_4887 = _T_4886 | _T_4760; // @[Mux.scala 27:72]
  wire  _T_4633 = ifu_ic_rw_int_addr_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire  _T_4761 = _T_4633 & way_status_out_13; // @[Mux.scala 27:72]
  wire  _T_4888 = _T_4887 | _T_4761; // @[Mux.scala 27:72]
  wire  _T_4634 = ifu_ic_rw_int_addr_ff == 7'he; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire  _T_4762 = _T_4634 & way_status_out_14; // @[Mux.scala 27:72]
  wire  _T_4889 = _T_4888 | _T_4762; // @[Mux.scala 27:72]
  wire  _T_4635 = ifu_ic_rw_int_addr_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire  _T_4763 = _T_4635 & way_status_out_15; // @[Mux.scala 27:72]
  wire  _T_4890 = _T_4889 | _T_4763; // @[Mux.scala 27:72]
  wire  _T_4636 = ifu_ic_rw_int_addr_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire  _T_4764 = _T_4636 & way_status_out_16; // @[Mux.scala 27:72]
  wire  _T_4891 = _T_4890 | _T_4764; // @[Mux.scala 27:72]
  wire  _T_4637 = ifu_ic_rw_int_addr_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire  _T_4765 = _T_4637 & way_status_out_17; // @[Mux.scala 27:72]
  wire  _T_4892 = _T_4891 | _T_4765; // @[Mux.scala 27:72]
  wire  _T_4638 = ifu_ic_rw_int_addr_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire  _T_4766 = _T_4638 & way_status_out_18; // @[Mux.scala 27:72]
  wire  _T_4893 = _T_4892 | _T_4766; // @[Mux.scala 27:72]
  wire  _T_4639 = ifu_ic_rw_int_addr_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire  _T_4767 = _T_4639 & way_status_out_19; // @[Mux.scala 27:72]
  wire  _T_4894 = _T_4893 | _T_4767; // @[Mux.scala 27:72]
  wire  _T_4640 = ifu_ic_rw_int_addr_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire  _T_4768 = _T_4640 & way_status_out_20; // @[Mux.scala 27:72]
  wire  _T_4895 = _T_4894 | _T_4768; // @[Mux.scala 27:72]
  wire  _T_4641 = ifu_ic_rw_int_addr_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire  _T_4769 = _T_4641 & way_status_out_21; // @[Mux.scala 27:72]
  wire  _T_4896 = _T_4895 | _T_4769; // @[Mux.scala 27:72]
  wire  _T_4642 = ifu_ic_rw_int_addr_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire  _T_4770 = _T_4642 & way_status_out_22; // @[Mux.scala 27:72]
  wire  _T_4897 = _T_4896 | _T_4770; // @[Mux.scala 27:72]
  wire  _T_4643 = ifu_ic_rw_int_addr_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire  _T_4771 = _T_4643 & way_status_out_23; // @[Mux.scala 27:72]
  wire  _T_4898 = _T_4897 | _T_4771; // @[Mux.scala 27:72]
  wire  _T_4644 = ifu_ic_rw_int_addr_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire  _T_4772 = _T_4644 & way_status_out_24; // @[Mux.scala 27:72]
  wire  _T_4899 = _T_4898 | _T_4772; // @[Mux.scala 27:72]
  wire  _T_4645 = ifu_ic_rw_int_addr_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire  _T_4773 = _T_4645 & way_status_out_25; // @[Mux.scala 27:72]
  wire  _T_4900 = _T_4899 | _T_4773; // @[Mux.scala 27:72]
  wire  _T_4646 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire  _T_4774 = _T_4646 & way_status_out_26; // @[Mux.scala 27:72]
  wire  _T_4901 = _T_4900 | _T_4774; // @[Mux.scala 27:72]
  wire  _T_4647 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire  _T_4775 = _T_4647 & way_status_out_27; // @[Mux.scala 27:72]
  wire  _T_4902 = _T_4901 | _T_4775; // @[Mux.scala 27:72]
  wire  _T_4648 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire  _T_4776 = _T_4648 & way_status_out_28; // @[Mux.scala 27:72]
  wire  _T_4903 = _T_4902 | _T_4776; // @[Mux.scala 27:72]
  wire  _T_4649 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire  _T_4777 = _T_4649 & way_status_out_29; // @[Mux.scala 27:72]
  wire  _T_4904 = _T_4903 | _T_4777; // @[Mux.scala 27:72]
  wire  _T_4650 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire  _T_4778 = _T_4650 & way_status_out_30; // @[Mux.scala 27:72]
  wire  _T_4905 = _T_4904 | _T_4778; // @[Mux.scala 27:72]
  wire  _T_4651 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire  _T_4779 = _T_4651 & way_status_out_31; // @[Mux.scala 27:72]
  wire  _T_4906 = _T_4905 | _T_4779; // @[Mux.scala 27:72]
  wire  _T_4652 = ifu_ic_rw_int_addr_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire  _T_4780 = _T_4652 & way_status_out_32; // @[Mux.scala 27:72]
  wire  _T_4907 = _T_4906 | _T_4780; // @[Mux.scala 27:72]
  wire  _T_4653 = ifu_ic_rw_int_addr_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire  _T_4781 = _T_4653 & way_status_out_33; // @[Mux.scala 27:72]
  wire  _T_4908 = _T_4907 | _T_4781; // @[Mux.scala 27:72]
  wire  _T_4654 = ifu_ic_rw_int_addr_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire  _T_4782 = _T_4654 & way_status_out_34; // @[Mux.scala 27:72]
  wire  _T_4909 = _T_4908 | _T_4782; // @[Mux.scala 27:72]
  wire  _T_4655 = ifu_ic_rw_int_addr_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire  _T_4783 = _T_4655 & way_status_out_35; // @[Mux.scala 27:72]
  wire  _T_4910 = _T_4909 | _T_4783; // @[Mux.scala 27:72]
  wire  _T_4656 = ifu_ic_rw_int_addr_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire  _T_4784 = _T_4656 & way_status_out_36; // @[Mux.scala 27:72]
  wire  _T_4911 = _T_4910 | _T_4784; // @[Mux.scala 27:72]
  wire  _T_4657 = ifu_ic_rw_int_addr_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire  _T_4785 = _T_4657 & way_status_out_37; // @[Mux.scala 27:72]
  wire  _T_4912 = _T_4911 | _T_4785; // @[Mux.scala 27:72]
  wire  _T_4658 = ifu_ic_rw_int_addr_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire  _T_4786 = _T_4658 & way_status_out_38; // @[Mux.scala 27:72]
  wire  _T_4913 = _T_4912 | _T_4786; // @[Mux.scala 27:72]
  wire  _T_4659 = ifu_ic_rw_int_addr_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire  _T_4787 = _T_4659 & way_status_out_39; // @[Mux.scala 27:72]
  wire  _T_4914 = _T_4913 | _T_4787; // @[Mux.scala 27:72]
  wire  _T_4660 = ifu_ic_rw_int_addr_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire  _T_4788 = _T_4660 & way_status_out_40; // @[Mux.scala 27:72]
  wire  _T_4915 = _T_4914 | _T_4788; // @[Mux.scala 27:72]
  wire  _T_4661 = ifu_ic_rw_int_addr_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire  _T_4789 = _T_4661 & way_status_out_41; // @[Mux.scala 27:72]
  wire  _T_4916 = _T_4915 | _T_4789; // @[Mux.scala 27:72]
  wire  _T_4662 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire  _T_4790 = _T_4662 & way_status_out_42; // @[Mux.scala 27:72]
  wire  _T_4917 = _T_4916 | _T_4790; // @[Mux.scala 27:72]
  wire  _T_4663 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire  _T_4791 = _T_4663 & way_status_out_43; // @[Mux.scala 27:72]
  wire  _T_4918 = _T_4917 | _T_4791; // @[Mux.scala 27:72]
  wire  _T_4664 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire  _T_4792 = _T_4664 & way_status_out_44; // @[Mux.scala 27:72]
  wire  _T_4919 = _T_4918 | _T_4792; // @[Mux.scala 27:72]
  wire  _T_4665 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire  _T_4793 = _T_4665 & way_status_out_45; // @[Mux.scala 27:72]
  wire  _T_4920 = _T_4919 | _T_4793; // @[Mux.scala 27:72]
  wire  _T_4666 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire  _T_4794 = _T_4666 & way_status_out_46; // @[Mux.scala 27:72]
  wire  _T_4921 = _T_4920 | _T_4794; // @[Mux.scala 27:72]
  wire  _T_4667 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire  _T_4795 = _T_4667 & way_status_out_47; // @[Mux.scala 27:72]
  wire  _T_4922 = _T_4921 | _T_4795; // @[Mux.scala 27:72]
  wire  _T_4668 = ifu_ic_rw_int_addr_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire  _T_4796 = _T_4668 & way_status_out_48; // @[Mux.scala 27:72]
  wire  _T_4923 = _T_4922 | _T_4796; // @[Mux.scala 27:72]
  wire  _T_4669 = ifu_ic_rw_int_addr_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire  _T_4797 = _T_4669 & way_status_out_49; // @[Mux.scala 27:72]
  wire  _T_4924 = _T_4923 | _T_4797; // @[Mux.scala 27:72]
  wire  _T_4670 = ifu_ic_rw_int_addr_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire  _T_4798 = _T_4670 & way_status_out_50; // @[Mux.scala 27:72]
  wire  _T_4925 = _T_4924 | _T_4798; // @[Mux.scala 27:72]
  wire  _T_4671 = ifu_ic_rw_int_addr_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire  _T_4799 = _T_4671 & way_status_out_51; // @[Mux.scala 27:72]
  wire  _T_4926 = _T_4925 | _T_4799; // @[Mux.scala 27:72]
  wire  _T_4672 = ifu_ic_rw_int_addr_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire  _T_4800 = _T_4672 & way_status_out_52; // @[Mux.scala 27:72]
  wire  _T_4927 = _T_4926 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4673 = ifu_ic_rw_int_addr_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire  _T_4801 = _T_4673 & way_status_out_53; // @[Mux.scala 27:72]
  wire  _T_4928 = _T_4927 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4674 = ifu_ic_rw_int_addr_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire  _T_4802 = _T_4674 & way_status_out_54; // @[Mux.scala 27:72]
  wire  _T_4929 = _T_4928 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4675 = ifu_ic_rw_int_addr_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire  _T_4803 = _T_4675 & way_status_out_55; // @[Mux.scala 27:72]
  wire  _T_4930 = _T_4929 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4676 = ifu_ic_rw_int_addr_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire  _T_4804 = _T_4676 & way_status_out_56; // @[Mux.scala 27:72]
  wire  _T_4931 = _T_4930 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4677 = ifu_ic_rw_int_addr_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire  _T_4805 = _T_4677 & way_status_out_57; // @[Mux.scala 27:72]
  wire  _T_4932 = _T_4931 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4678 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire  _T_4806 = _T_4678 & way_status_out_58; // @[Mux.scala 27:72]
  wire  _T_4933 = _T_4932 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4679 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire  _T_4807 = _T_4679 & way_status_out_59; // @[Mux.scala 27:72]
  wire  _T_4934 = _T_4933 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4680 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire  _T_4808 = _T_4680 & way_status_out_60; // @[Mux.scala 27:72]
  wire  _T_4935 = _T_4934 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4681 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire  _T_4809 = _T_4681 & way_status_out_61; // @[Mux.scala 27:72]
  wire  _T_4936 = _T_4935 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4682 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire  _T_4810 = _T_4682 & way_status_out_62; // @[Mux.scala 27:72]
  wire  _T_4937 = _T_4936 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4683 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire  _T_4811 = _T_4683 & way_status_out_63; // @[Mux.scala 27:72]
  wire  _T_4938 = _T_4937 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4684 = ifu_ic_rw_int_addr_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire  _T_4812 = _T_4684 & way_status_out_64; // @[Mux.scala 27:72]
  wire  _T_4939 = _T_4938 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4685 = ifu_ic_rw_int_addr_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire  _T_4813 = _T_4685 & way_status_out_65; // @[Mux.scala 27:72]
  wire  _T_4940 = _T_4939 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4686 = ifu_ic_rw_int_addr_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire  _T_4814 = _T_4686 & way_status_out_66; // @[Mux.scala 27:72]
  wire  _T_4941 = _T_4940 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4687 = ifu_ic_rw_int_addr_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire  _T_4815 = _T_4687 & way_status_out_67; // @[Mux.scala 27:72]
  wire  _T_4942 = _T_4941 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4688 = ifu_ic_rw_int_addr_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire  _T_4816 = _T_4688 & way_status_out_68; // @[Mux.scala 27:72]
  wire  _T_4943 = _T_4942 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4689 = ifu_ic_rw_int_addr_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire  _T_4817 = _T_4689 & way_status_out_69; // @[Mux.scala 27:72]
  wire  _T_4944 = _T_4943 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4690 = ifu_ic_rw_int_addr_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire  _T_4818 = _T_4690 & way_status_out_70; // @[Mux.scala 27:72]
  wire  _T_4945 = _T_4944 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4691 = ifu_ic_rw_int_addr_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire  _T_4819 = _T_4691 & way_status_out_71; // @[Mux.scala 27:72]
  wire  _T_4946 = _T_4945 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4692 = ifu_ic_rw_int_addr_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire  _T_4820 = _T_4692 & way_status_out_72; // @[Mux.scala 27:72]
  wire  _T_4947 = _T_4946 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4693 = ifu_ic_rw_int_addr_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire  _T_4821 = _T_4693 & way_status_out_73; // @[Mux.scala 27:72]
  wire  _T_4948 = _T_4947 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4694 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire  _T_4822 = _T_4694 & way_status_out_74; // @[Mux.scala 27:72]
  wire  _T_4949 = _T_4948 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4695 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire  _T_4823 = _T_4695 & way_status_out_75; // @[Mux.scala 27:72]
  wire  _T_4950 = _T_4949 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4696 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire  _T_4824 = _T_4696 & way_status_out_76; // @[Mux.scala 27:72]
  wire  _T_4951 = _T_4950 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4697 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire  _T_4825 = _T_4697 & way_status_out_77; // @[Mux.scala 27:72]
  wire  _T_4952 = _T_4951 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4698 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire  _T_4826 = _T_4698 & way_status_out_78; // @[Mux.scala 27:72]
  wire  _T_4953 = _T_4952 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4699 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire  _T_4827 = _T_4699 & way_status_out_79; // @[Mux.scala 27:72]
  wire  _T_4954 = _T_4953 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4700 = ifu_ic_rw_int_addr_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire  _T_4828 = _T_4700 & way_status_out_80; // @[Mux.scala 27:72]
  wire  _T_4955 = _T_4954 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4701 = ifu_ic_rw_int_addr_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire  _T_4829 = _T_4701 & way_status_out_81; // @[Mux.scala 27:72]
  wire  _T_4956 = _T_4955 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4702 = ifu_ic_rw_int_addr_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire  _T_4830 = _T_4702 & way_status_out_82; // @[Mux.scala 27:72]
  wire  _T_4957 = _T_4956 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4703 = ifu_ic_rw_int_addr_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire  _T_4831 = _T_4703 & way_status_out_83; // @[Mux.scala 27:72]
  wire  _T_4958 = _T_4957 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4704 = ifu_ic_rw_int_addr_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire  _T_4832 = _T_4704 & way_status_out_84; // @[Mux.scala 27:72]
  wire  _T_4959 = _T_4958 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4705 = ifu_ic_rw_int_addr_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire  _T_4833 = _T_4705 & way_status_out_85; // @[Mux.scala 27:72]
  wire  _T_4960 = _T_4959 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4706 = ifu_ic_rw_int_addr_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire  _T_4834 = _T_4706 & way_status_out_86; // @[Mux.scala 27:72]
  wire  _T_4961 = _T_4960 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4707 = ifu_ic_rw_int_addr_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire  _T_4835 = _T_4707 & way_status_out_87; // @[Mux.scala 27:72]
  wire  _T_4962 = _T_4961 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4708 = ifu_ic_rw_int_addr_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire  _T_4836 = _T_4708 & way_status_out_88; // @[Mux.scala 27:72]
  wire  _T_4963 = _T_4962 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4709 = ifu_ic_rw_int_addr_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire  _T_4837 = _T_4709 & way_status_out_89; // @[Mux.scala 27:72]
  wire  _T_4964 = _T_4963 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4710 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire  _T_4838 = _T_4710 & way_status_out_90; // @[Mux.scala 27:72]
  wire  _T_4965 = _T_4964 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4711 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire  _T_4839 = _T_4711 & way_status_out_91; // @[Mux.scala 27:72]
  wire  _T_4966 = _T_4965 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4712 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire  _T_4840 = _T_4712 & way_status_out_92; // @[Mux.scala 27:72]
  wire  _T_4967 = _T_4966 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4713 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire  _T_4841 = _T_4713 & way_status_out_93; // @[Mux.scala 27:72]
  wire  _T_4968 = _T_4967 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4714 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire  _T_4842 = _T_4714 & way_status_out_94; // @[Mux.scala 27:72]
  wire  _T_4969 = _T_4968 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4715 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire  _T_4843 = _T_4715 & way_status_out_95; // @[Mux.scala 27:72]
  wire  _T_4970 = _T_4969 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4716 = ifu_ic_rw_int_addr_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire  _T_4844 = _T_4716 & way_status_out_96; // @[Mux.scala 27:72]
  wire  _T_4971 = _T_4970 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4717 = ifu_ic_rw_int_addr_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire  _T_4845 = _T_4717 & way_status_out_97; // @[Mux.scala 27:72]
  wire  _T_4972 = _T_4971 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4718 = ifu_ic_rw_int_addr_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire  _T_4846 = _T_4718 & way_status_out_98; // @[Mux.scala 27:72]
  wire  _T_4973 = _T_4972 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4719 = ifu_ic_rw_int_addr_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire  _T_4847 = _T_4719 & way_status_out_99; // @[Mux.scala 27:72]
  wire  _T_4974 = _T_4973 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4720 = ifu_ic_rw_int_addr_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire  _T_4848 = _T_4720 & way_status_out_100; // @[Mux.scala 27:72]
  wire  _T_4975 = _T_4974 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4721 = ifu_ic_rw_int_addr_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire  _T_4849 = _T_4721 & way_status_out_101; // @[Mux.scala 27:72]
  wire  _T_4976 = _T_4975 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4722 = ifu_ic_rw_int_addr_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire  _T_4850 = _T_4722 & way_status_out_102; // @[Mux.scala 27:72]
  wire  _T_4977 = _T_4976 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4723 = ifu_ic_rw_int_addr_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire  _T_4851 = _T_4723 & way_status_out_103; // @[Mux.scala 27:72]
  wire  _T_4978 = _T_4977 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4724 = ifu_ic_rw_int_addr_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire  _T_4852 = _T_4724 & way_status_out_104; // @[Mux.scala 27:72]
  wire  _T_4979 = _T_4978 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4725 = ifu_ic_rw_int_addr_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire  _T_4853 = _T_4725 & way_status_out_105; // @[Mux.scala 27:72]
  wire  _T_4980 = _T_4979 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4726 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire  _T_4854 = _T_4726 & way_status_out_106; // @[Mux.scala 27:72]
  wire  _T_4981 = _T_4980 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4727 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire  _T_4855 = _T_4727 & way_status_out_107; // @[Mux.scala 27:72]
  wire  _T_4982 = _T_4981 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4728 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire  _T_4856 = _T_4728 & way_status_out_108; // @[Mux.scala 27:72]
  wire  _T_4983 = _T_4982 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4729 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire  _T_4857 = _T_4729 & way_status_out_109; // @[Mux.scala 27:72]
  wire  _T_4984 = _T_4983 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4730 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire  _T_4858 = _T_4730 & way_status_out_110; // @[Mux.scala 27:72]
  wire  _T_4985 = _T_4984 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4731 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire  _T_4859 = _T_4731 & way_status_out_111; // @[Mux.scala 27:72]
  wire  _T_4986 = _T_4985 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4732 = ifu_ic_rw_int_addr_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire  _T_4860 = _T_4732 & way_status_out_112; // @[Mux.scala 27:72]
  wire  _T_4987 = _T_4986 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4733 = ifu_ic_rw_int_addr_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire  _T_4861 = _T_4733 & way_status_out_113; // @[Mux.scala 27:72]
  wire  _T_4988 = _T_4987 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4734 = ifu_ic_rw_int_addr_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire  _T_4862 = _T_4734 & way_status_out_114; // @[Mux.scala 27:72]
  wire  _T_4989 = _T_4988 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4735 = ifu_ic_rw_int_addr_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire  _T_4863 = _T_4735 & way_status_out_115; // @[Mux.scala 27:72]
  wire  _T_4990 = _T_4989 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4736 = ifu_ic_rw_int_addr_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire  _T_4864 = _T_4736 & way_status_out_116; // @[Mux.scala 27:72]
  wire  _T_4991 = _T_4990 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4737 = ifu_ic_rw_int_addr_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire  _T_4865 = _T_4737 & way_status_out_117; // @[Mux.scala 27:72]
  wire  _T_4992 = _T_4991 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4738 = ifu_ic_rw_int_addr_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire  _T_4866 = _T_4738 & way_status_out_118; // @[Mux.scala 27:72]
  wire  _T_4993 = _T_4992 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4739 = ifu_ic_rw_int_addr_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire  _T_4867 = _T_4739 & way_status_out_119; // @[Mux.scala 27:72]
  wire  _T_4994 = _T_4993 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4740 = ifu_ic_rw_int_addr_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire  _T_4868 = _T_4740 & way_status_out_120; // @[Mux.scala 27:72]
  wire  _T_4995 = _T_4994 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4741 = ifu_ic_rw_int_addr_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire  _T_4869 = _T_4741 & way_status_out_121; // @[Mux.scala 27:72]
  wire  _T_4996 = _T_4995 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4742 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire  _T_4870 = _T_4742 & way_status_out_122; // @[Mux.scala 27:72]
  wire  _T_4997 = _T_4996 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4743 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire  _T_4871 = _T_4743 & way_status_out_123; // @[Mux.scala 27:72]
  wire  _T_4998 = _T_4997 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4744 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire  _T_4872 = _T_4744 & way_status_out_124; // @[Mux.scala 27:72]
  wire  _T_4999 = _T_4998 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4745 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire  _T_4873 = _T_4745 & way_status_out_125; // @[Mux.scala 27:72]
  wire  _T_5000 = _T_4999 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4746 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire  _T_4874 = _T_4746 & way_status_out_126; // @[Mux.scala 27:72]
  wire  _T_5001 = _T_5000 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_4747 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 733:80]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire  _T_4875 = _T_4747 & way_status_out_127; // @[Mux.scala 27:72]
  wire  way_status = _T_5001 | _T_4875; // @[Mux.scala 27:72]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 263:96]
  wire [1:0] _T_197 = _T_195 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_198 = _T_197 & io_ic_tag_valid; // @[el2_ifu_mem_ctl.scala 263:113]
  reg [1:0] tagv_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 269:58]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 265:67]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:54]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[el2_ifu_mem_ctl.scala 583:46]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 272:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 277:59]
  wire  _T_214 = _T_212 | _T_2219; // @[el2_ifu_mem_ctl.scala 277:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 277:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 283:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 283:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 283:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 290:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 290:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 290:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 291:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 291:32]
  wire  _T_274 = imb_ff[11:5] == imb_scnd_ff[11:5]; // @[el2_ifu_mem_ctl.scala 294:79]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 294:135]
  reg [1:0] ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 581:51]
  wire  _T_2644 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 626:48]
  wire  _T_2645 = _T_2644 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 626:52]
  wire  bus_ifu_wr_data_error_ff = _T_2645 & miss_pending; // @[el2_ifu_mem_ctl.scala 626:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 368:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 367:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 294:153]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 294:151]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 297:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 297:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 298:24]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 318:59]
  wire  _T_9705 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 789:31]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 319:53]
  wire  _T_9707 = _T_9705 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 789:49]
  wire  _T_9709 = _T_9707 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 789:65]
  wire  _T_9711 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 789:84]
  wire  replace_way_mb_any_0 = _T_9709 | _T_9711; // @[el2_ifu_mem_ctl.scala 789:82]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9714 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 790:48]
  wire  _T_9716 = _T_9714 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 790:64]
  wire  _T_9718 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 790:83]
  wire  _T_9720 = _T_9718 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 790:98]
  wire  replace_way_mb_any_1 = _T_9716 | _T_9720; // @[el2_ifu_mem_ctl.scala 790:81]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 302:110]
  wire [1:0] _T_290 = tagv_mb_scnd_ff | _T_289; // @[el2_ifu_mem_ctl.scala 302:62]
  wire [1:0] _T_295 = io_ic_tag_valid & _T_197; // @[el2_ifu_mem_ctl.scala 303:58]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 306:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 306:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 307:48]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 306:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 306:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 308:62]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 317:48]
  wire  _T_309 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 316:57]
  wire  _T_315 = _T_2234 & flush_final_f; // @[el2_ifu_mem_ctl.scala 321:87]
  wire  _T_316 = ~_T_315; // @[el2_ifu_mem_ctl.scala 321:55]
  wire  _T_317 = io_ifc_fetch_req_bf & _T_316; // @[el2_ifu_mem_ctl.scala 321:53]
  wire  _T_2226 = ~_T_2221; // @[el2_ifu_mem_ctl.scala 459:46]
  wire  _T_2227 = _T_2219 & _T_2226; // @[el2_ifu_mem_ctl.scala 459:44]
  wire  stream_miss_f = _T_2227 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 459:84]
  wire  _T_318 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 321:106]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 327:68]
  reg [2:0] bus_rd_addr_count; // @[el2_ifu_mem_ctl.scala 608:55]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_325 = _T_239 | _T_2219; // @[el2_ifu_mem_ctl.scala 329:55]
  wire  _T_328 = _T_325 & _T_56; // @[el2_ifu_mem_ctl.scala 329:82]
  wire  _T_2240 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 464:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2240}; // @[Cat.scala 29:58]
  wire  _T_2241 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 465:81]
  wire  _T_2265 = _T_2241 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2244 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 465:81]
  wire  _T_2266 = _T_2244 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2273 = _T_2265 | _T_2266; // @[Mux.scala 27:72]
  wire  _T_2247 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 465:81]
  wire  _T_2267 = _T_2247 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2274 = _T_2273 | _T_2267; // @[Mux.scala 27:72]
  wire  _T_2250 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 465:81]
  wire  _T_2268 = _T_2250 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2275 = _T_2274 | _T_2268; // @[Mux.scala 27:72]
  wire  _T_2253 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 465:81]
  wire  _T_2269 = _T_2253 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2276 = _T_2275 | _T_2269; // @[Mux.scala 27:72]
  wire  _T_2256 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 465:81]
  wire  _T_2270 = _T_2256 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2277 = _T_2276 | _T_2270; // @[Mux.scala 27:72]
  wire  _T_2259 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 465:81]
  wire  _T_2271 = _T_2259 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2278 = _T_2277 | _T_2271; // @[Mux.scala 27:72]
  wire  _T_2262 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 465:81]
  wire  _T_2272 = _T_2262 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2278 | _T_2272; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 466:46]
  wire  _T_332 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 333:35]
  wire  _T_334 = _T_332 & _T_17; // @[el2_ifu_mem_ctl.scala 333:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 623:61]
  wire  _T_2638 = ic_act_miss_f_delayed & _T_2235; // @[el2_ifu_mem_ctl.scala 624:53]
  wire  reset_tag_valid_for_miss = _T_2638 & _T_17; // @[el2_ifu_mem_ctl.scala 624:84]
  wire  sel_mb_addr = _T_334 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 333:79]
  wire [30:0] _T_338 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_339 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 335:5]
  wire [30:0] _T_340 = sel_mb_addr ? _T_338 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_341 = _T_339 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_340 | _T_341; // @[Mux.scala 27:72]
  wire  _T_346 = _T_334 & last_beat; // @[el2_ifu_mem_ctl.scala 337:84]
  wire  _T_2632 = ~_T_2644; // @[el2_ifu_mem_ctl.scala 621:84]
  wire  _T_2633 = _T_100 & _T_2632; // @[el2_ifu_mem_ctl.scala 621:82]
  wire  bus_ifu_wr_en_ff_q = _T_2633 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 621:108]
  wire  sel_mb_status_addr = _T_346 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 337:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_338 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 338:31]
  reg [63:0] ifu_bus_rdata_ff; // @[el2_ifu_mem_ctl.scala 582:48]
  wire [6:0] _T_569 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 416:13]
  wire  _T_570 = ^_T_569; // @[el2_lib.scala 416:20]
  wire [6:0] _T_576 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_583 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 416:30]
  wire [14:0] _T_584 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_576}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_591 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 416:30]
  wire [30:0] _T_600 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_591,_T_584}; // @[el2_lib.scala 416:30]
  wire  _T_601 = ^_T_600; // @[el2_lib.scala 416:37]
  wire [6:0] _T_607 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 416:47]
  wire [14:0] _T_615 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_607}; // @[el2_lib.scala 416:47]
  wire [30:0] _T_631 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_591,_T_615}; // @[el2_lib.scala 416:47]
  wire  _T_632 = ^_T_631; // @[el2_lib.scala 416:54]
  wire [6:0] _T_638 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 416:64]
  wire [14:0] _T_646 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_638}; // @[el2_lib.scala 416:64]
  wire [30:0] _T_662 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_583,_T_646}; // @[el2_lib.scala 416:64]
  wire  _T_663 = ^_T_662; // @[el2_lib.scala 416:71]
  wire [7:0] _T_670 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 416:81]
  wire [16:0] _T_679 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_670}; // @[el2_lib.scala 416:81]
  wire [8:0] _T_687 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 416:81]
  wire [17:0] _T_696 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_687}; // @[el2_lib.scala 416:81]
  wire [34:0] _T_697 = {_T_696,_T_679}; // @[el2_lib.scala 416:81]
  wire  _T_698 = ^_T_697; // @[el2_lib.scala 416:88]
  wire [7:0] _T_705 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 416:98]
  wire [16:0] _T_714 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_705}; // @[el2_lib.scala 416:98]
  wire [8:0] _T_722 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 416:98]
  wire [17:0] _T_731 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_722}; // @[el2_lib.scala 416:98]
  wire [34:0] _T_732 = {_T_731,_T_714}; // @[el2_lib.scala 416:98]
  wire  _T_733 = ^_T_732; // @[el2_lib.scala 416:105]
  wire [7:0] _T_740 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 416:115]
  wire [16:0] _T_749 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_740}; // @[el2_lib.scala 416:115]
  wire [8:0] _T_757 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 416:115]
  wire [17:0] _T_766 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_757}; // @[el2_lib.scala 416:115]
  wire [34:0] _T_767 = {_T_766,_T_749}; // @[el2_lib.scala 416:115]
  wire  _T_768 = ^_T_767; // @[el2_lib.scala 416:122]
  wire [3:0] _T_2281 = {ifu_bus_rid_ff[2:1],_T_2240,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2282 = _T_2281 == 4'h0; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_0; // @[el2_ifu_mem_ctl.scala 402:67]
  wire [31:0] _T_2329 = _T_2282 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2285 = _T_2281 == 4'h1; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_1; // @[el2_ifu_mem_ctl.scala 403:69]
  wire [31:0] _T_2330 = _T_2285 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2345 = _T_2329 | _T_2330; // @[Mux.scala 27:72]
  wire  _T_2288 = _T_2281 == 4'h2; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_2; // @[el2_ifu_mem_ctl.scala 402:67]
  wire [31:0] _T_2331 = _T_2288 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2346 = _T_2345 | _T_2331; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2281 == 4'h3; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_3; // @[el2_ifu_mem_ctl.scala 403:69]
  wire [31:0] _T_2332 = _T_2291 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2347 = _T_2346 | _T_2332; // @[Mux.scala 27:72]
  wire  _T_2294 = _T_2281 == 4'h4; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_4; // @[el2_ifu_mem_ctl.scala 402:67]
  wire [31:0] _T_2333 = _T_2294 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2348 = _T_2347 | _T_2333; // @[Mux.scala 27:72]
  wire  _T_2297 = _T_2281 == 4'h5; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_5; // @[el2_ifu_mem_ctl.scala 403:69]
  wire [31:0] _T_2334 = _T_2297 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2349 = _T_2348 | _T_2334; // @[Mux.scala 27:72]
  wire  _T_2300 = _T_2281 == 4'h6; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_6; // @[el2_ifu_mem_ctl.scala 402:67]
  wire [31:0] _T_2335 = _T_2300 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2350 = _T_2349 | _T_2335; // @[Mux.scala 27:72]
  wire  _T_2303 = _T_2281 == 4'h7; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_7; // @[el2_ifu_mem_ctl.scala 403:69]
  wire [31:0] _T_2336 = _T_2303 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2351 = _T_2350 | _T_2336; // @[Mux.scala 27:72]
  wire  _T_2306 = _T_2281 == 4'h8; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_8; // @[el2_ifu_mem_ctl.scala 402:67]
  wire [31:0] _T_2337 = _T_2306 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2352 = _T_2351 | _T_2337; // @[Mux.scala 27:72]
  wire  _T_2309 = _T_2281 == 4'h9; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_9; // @[el2_ifu_mem_ctl.scala 403:69]
  wire [31:0] _T_2338 = _T_2309 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2353 = _T_2352 | _T_2338; // @[Mux.scala 27:72]
  wire  _T_2312 = _T_2281 == 4'ha; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_10; // @[el2_ifu_mem_ctl.scala 402:67]
  wire [31:0] _T_2339 = _T_2312 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2354 = _T_2353 | _T_2339; // @[Mux.scala 27:72]
  wire  _T_2315 = _T_2281 == 4'hb; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_11; // @[el2_ifu_mem_ctl.scala 403:69]
  wire [31:0] _T_2340 = _T_2315 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2355 = _T_2354 | _T_2340; // @[Mux.scala 27:72]
  wire  _T_2318 = _T_2281 == 4'hc; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_12; // @[el2_ifu_mem_ctl.scala 402:67]
  wire [31:0] _T_2341 = _T_2318 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2356 = _T_2355 | _T_2341; // @[Mux.scala 27:72]
  wire  _T_2321 = _T_2281 == 4'hd; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_13; // @[el2_ifu_mem_ctl.scala 403:69]
  wire [31:0] _T_2342 = _T_2321 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2357 = _T_2356 | _T_2342; // @[Mux.scala 27:72]
  wire  _T_2324 = _T_2281 == 4'he; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_14; // @[el2_ifu_mem_ctl.scala 402:67]
  wire [31:0] _T_2343 = _T_2324 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2358 = _T_2357 | _T_2343; // @[Mux.scala 27:72]
  wire  _T_2327 = _T_2281 == 4'hf; // @[el2_ifu_mem_ctl.scala 467:89]
  reg [31:0] ic_miss_buff_data_15; // @[el2_ifu_mem_ctl.scala 403:69]
  wire [31:0] _T_2344 = _T_2327 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2359 = _T_2358 | _T_2344; // @[Mux.scala 27:72]
  wire [3:0] _T_2361 = {ifu_bus_rid_ff[2:1],_T_2240,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2362 = _T_2361 == 4'h0; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2409 = _T_2362 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2365 = _T_2361 == 4'h1; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2410 = _T_2365 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2425 = _T_2409 | _T_2410; // @[Mux.scala 27:72]
  wire  _T_2368 = _T_2361 == 4'h2; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2411 = _T_2368 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2426 = _T_2425 | _T_2411; // @[Mux.scala 27:72]
  wire  _T_2371 = _T_2361 == 4'h3; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2412 = _T_2371 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2427 = _T_2426 | _T_2412; // @[Mux.scala 27:72]
  wire  _T_2374 = _T_2361 == 4'h4; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2413 = _T_2374 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2428 = _T_2427 | _T_2413; // @[Mux.scala 27:72]
  wire  _T_2377 = _T_2361 == 4'h5; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2414 = _T_2377 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2429 = _T_2428 | _T_2414; // @[Mux.scala 27:72]
  wire  _T_2380 = _T_2361 == 4'h6; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2415 = _T_2380 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2430 = _T_2429 | _T_2415; // @[Mux.scala 27:72]
  wire  _T_2383 = _T_2361 == 4'h7; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2416 = _T_2383 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2431 = _T_2430 | _T_2416; // @[Mux.scala 27:72]
  wire  _T_2386 = _T_2361 == 4'h8; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2417 = _T_2386 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2432 = _T_2431 | _T_2417; // @[Mux.scala 27:72]
  wire  _T_2389 = _T_2361 == 4'h9; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2418 = _T_2389 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2433 = _T_2432 | _T_2418; // @[Mux.scala 27:72]
  wire  _T_2392 = _T_2361 == 4'ha; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2419 = _T_2392 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2434 = _T_2433 | _T_2419; // @[Mux.scala 27:72]
  wire  _T_2395 = _T_2361 == 4'hb; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2420 = _T_2395 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2435 = _T_2434 | _T_2420; // @[Mux.scala 27:72]
  wire  _T_2398 = _T_2361 == 4'hc; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2421 = _T_2398 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2436 = _T_2435 | _T_2421; // @[Mux.scala 27:72]
  wire  _T_2401 = _T_2361 == 4'hd; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2422 = _T_2401 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2437 = _T_2436 | _T_2422; // @[Mux.scala 27:72]
  wire  _T_2404 = _T_2361 == 4'he; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2423 = _T_2404 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2438 = _T_2437 | _T_2423; // @[Mux.scala 27:72]
  wire  _T_2407 = _T_2361 == 4'hf; // @[el2_ifu_mem_ctl.scala 468:66]
  wire [31:0] _T_2424 = _T_2407 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2439 = _T_2438 | _T_2424; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2359,_T_2439}; // @[Cat.scala 29:58]
  wire [6:0] _T_991 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 416:13]
  wire  _T_992 = ^_T_991; // @[el2_lib.scala 416:20]
  wire [6:0] _T_998 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_1005 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 416:30]
  wire [14:0] _T_1006 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_998}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_1013 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 416:30]
  wire [30:0] _T_1022 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1013,_T_1006}; // @[el2_lib.scala 416:30]
  wire  _T_1023 = ^_T_1022; // @[el2_lib.scala 416:37]
  wire [6:0] _T_1029 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 416:47]
  wire [14:0] _T_1037 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1029}; // @[el2_lib.scala 416:47]
  wire [30:0] _T_1053 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1013,_T_1037}; // @[el2_lib.scala 416:47]
  wire  _T_1054 = ^_T_1053; // @[el2_lib.scala 416:54]
  wire [6:0] _T_1060 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 416:64]
  wire [14:0] _T_1068 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1060}; // @[el2_lib.scala 416:64]
  wire [30:0] _T_1084 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1005,_T_1068}; // @[el2_lib.scala 416:64]
  wire  _T_1085 = ^_T_1084; // @[el2_lib.scala 416:71]
  wire [7:0] _T_1092 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 416:81]
  wire [16:0] _T_1101 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1092}; // @[el2_lib.scala 416:81]
  wire [8:0] _T_1109 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 416:81]
  wire [17:0] _T_1118 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1109}; // @[el2_lib.scala 416:81]
  wire [34:0] _T_1119 = {_T_1118,_T_1101}; // @[el2_lib.scala 416:81]
  wire  _T_1120 = ^_T_1119; // @[el2_lib.scala 416:88]
  wire [7:0] _T_1127 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 416:98]
  wire [16:0] _T_1136 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1127}; // @[el2_lib.scala 416:98]
  wire [8:0] _T_1144 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 416:98]
  wire [17:0] _T_1153 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1144}; // @[el2_lib.scala 416:98]
  wire [34:0] _T_1154 = {_T_1153,_T_1136}; // @[el2_lib.scala 416:98]
  wire  _T_1155 = ^_T_1154; // @[el2_lib.scala 416:105]
  wire [7:0] _T_1162 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 416:115]
  wire [16:0] _T_1171 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1162}; // @[el2_lib.scala 416:115]
  wire [8:0] _T_1179 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 416:115]
  wire [17:0] _T_1188 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1179}; // @[el2_lib.scala 416:115]
  wire [34:0] _T_1189 = {_T_1188,_T_1171}; // @[el2_lib.scala 416:115]
  wire  _T_1190 = ^_T_1189; // @[el2_lib.scala 416:122]
  wire [70:0] _T_1235 = {_T_570,_T_601,_T_632,_T_663,_T_698,_T_733,_T_768,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1234 = {_T_992,_T_1023,_T_1054,_T_1085,_T_1120,_T_1155,_T_1190,_T_2359,_T_2439}; // @[Cat.scala 29:58]
  wire [141:0] _T_1236 = {_T_570,_T_601,_T_632,_T_663,_T_698,_T_733,_T_768,ifu_bus_rdata_ff,_T_1234}; // @[Cat.scala 29:58]
  wire [141:0] _T_1239 = {_T_992,_T_1023,_T_1054,_T_1085,_T_1120,_T_1155,_T_1190,_T_2359,_T_2439,_T_1235}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1236 : _T_1239; // @[el2_ifu_mem_ctl.scala 359:28]
  wire  _T_1198 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 349:56]
  wire  _T_1199 = _T_1198 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 349:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 414:28]
  wire  _T_1399 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 416:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 619:35]
  wire  _T_1284 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 398:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 398:73]
  wire  _T_1325 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 405:118]
  wire  _T_1326 = ic_miss_buff_data_valid[0] & _T_1325; // @[el2_ifu_mem_ctl.scala 405:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1326; // @[el2_ifu_mem_ctl.scala 405:88]
  wire  _T_1422 = _T_1399 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1402 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 416:114]
  wire  _T_1285 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 398:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1285; // @[el2_ifu_mem_ctl.scala 398:73]
  wire  _T_1329 = ic_miss_buff_data_valid[1] & _T_1325; // @[el2_ifu_mem_ctl.scala 405:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1329; // @[el2_ifu_mem_ctl.scala 405:88]
  wire  _T_1423 = _T_1402 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1430 = _T_1422 | _T_1423; // @[Mux.scala 27:72]
  wire  _T_1405 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 416:114]
  wire  _T_1286 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 398:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1286; // @[el2_ifu_mem_ctl.scala 398:73]
  wire  _T_1332 = ic_miss_buff_data_valid[2] & _T_1325; // @[el2_ifu_mem_ctl.scala 405:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1332; // @[el2_ifu_mem_ctl.scala 405:88]
  wire  _T_1424 = _T_1405 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1431 = _T_1430 | _T_1424; // @[Mux.scala 27:72]
  wire  _T_1408 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 416:114]
  wire  _T_1287 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 398:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 398:73]
  wire  _T_1335 = ic_miss_buff_data_valid[3] & _T_1325; // @[el2_ifu_mem_ctl.scala 405:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1335; // @[el2_ifu_mem_ctl.scala 405:88]
  wire  _T_1425 = _T_1408 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1432 = _T_1431 | _T_1425; // @[Mux.scala 27:72]
  wire  _T_1411 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 416:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 398:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 398:73]
  wire  _T_1338 = ic_miss_buff_data_valid[4] & _T_1325; // @[el2_ifu_mem_ctl.scala 405:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1338; // @[el2_ifu_mem_ctl.scala 405:88]
  wire  _T_1426 = _T_1411 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1433 = _T_1432 | _T_1426; // @[Mux.scala 27:72]
  wire  _T_1414 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 416:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 398:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 398:73]
  wire  _T_1341 = ic_miss_buff_data_valid[5] & _T_1325; // @[el2_ifu_mem_ctl.scala 405:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1341; // @[el2_ifu_mem_ctl.scala 405:88]
  wire  _T_1427 = _T_1414 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1434 = _T_1433 | _T_1427; // @[Mux.scala 27:72]
  wire  _T_1417 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 416:114]
  wire  _T_1290 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 398:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1290; // @[el2_ifu_mem_ctl.scala 398:73]
  wire  _T_1344 = ic_miss_buff_data_valid[6] & _T_1325; // @[el2_ifu_mem_ctl.scala 405:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1344; // @[el2_ifu_mem_ctl.scala 405:88]
  wire  _T_1428 = _T_1417 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1435 = _T_1434 | _T_1428; // @[Mux.scala 27:72]
  wire  _T_1420 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 416:114]
  wire  _T_1291 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 398:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1291; // @[el2_ifu_mem_ctl.scala 398:73]
  wire  _T_1347 = ic_miss_buff_data_valid[7] & _T_1325; // @[el2_ifu_mem_ctl.scala 405:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1347; // @[el2_ifu_mem_ctl.scala 405:88]
  wire  _T_1429 = _T_1420 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1435 | _T_1429; // @[Mux.scala 27:72]
  wire  _T_1438 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 417:58]
  wire  _T_1439 = bypass_valid_value_check & _T_1438; // @[el2_ifu_mem_ctl.scala 417:56]
  wire  _T_1441 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 417:77]
  wire  _T_1442 = _T_1439 & _T_1441; // @[el2_ifu_mem_ctl.scala 417:75]
  wire  _T_1447 = _T_1439 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 418:50]
  wire  _T_1448 = _T_1442 | _T_1447; // @[el2_ifu_mem_ctl.scala 417:95]
  wire  _T_1450 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 419:31]
  wire  _T_1453 = _T_1450 & _T_1441; // @[el2_ifu_mem_ctl.scala 419:49]
  wire  _T_1454 = _T_1448 | _T_1453; // @[el2_ifu_mem_ctl.scala 418:69]
  wire  _T_1458 = _T_1450 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 420:49]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 415:70]
  wire  _T_1459 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 420:130]
  wire  _T_1475 = _T_1459 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1461 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 420:130]
  wire  _T_1476 = _T_1461 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1483 = _T_1475 | _T_1476; // @[Mux.scala 27:72]
  wire  _T_1463 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 420:130]
  wire  _T_1477 = _T_1463 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1484 = _T_1483 | _T_1477; // @[Mux.scala 27:72]
  wire  _T_1465 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 420:130]
  wire  _T_1478 = _T_1465 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1485 = _T_1484 | _T_1478; // @[Mux.scala 27:72]
  wire  _T_1467 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 420:130]
  wire  _T_1479 = _T_1467 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1486 = _T_1485 | _T_1479; // @[Mux.scala 27:72]
  wire  _T_1469 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 420:130]
  wire  _T_1480 = _T_1469 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1487 = _T_1486 | _T_1480; // @[Mux.scala 27:72]
  wire  _T_1471 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 420:130]
  wire  _T_1481 = _T_1471 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1488 = _T_1487 | _T_1481; // @[Mux.scala 27:72]
  wire  _T_1473 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 420:130]
  wire  _T_1482 = _T_1473 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1489 = _T_1488 | _T_1482; // @[Mux.scala 27:72]
  wire  _T_1491 = _T_1458 & _T_1489; // @[el2_ifu_mem_ctl.scala 420:67]
  wire  _T_1492 = _T_1454 | _T_1491; // @[el2_ifu_mem_ctl.scala 419:69]
  wire [4:0] _GEN_446 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 421:70]
  wire  _T_1495 = _GEN_446 == 5'h1f; // @[el2_ifu_mem_ctl.scala 421:70]
  wire  _T_1496 = bypass_valid_value_check & _T_1495; // @[el2_ifu_mem_ctl.scala 421:31]
  wire  bypass_data_ready_in = _T_1492 | _T_1496; // @[el2_ifu_mem_ctl.scala 420:179]
  wire  _T_1497 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 425:53]
  wire  _T_1498 = _T_1497 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 425:73]
  wire  _T_1500 = _T_1498 & _T_319; // @[el2_ifu_mem_ctl.scala 425:96]
  wire  _T_1502 = _T_1500 & _T_58; // @[el2_ifu_mem_ctl.scala 425:118]
  wire  _T_1504 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 426:47]
  wire  _T_1506 = _T_1504 & _T_319; // @[el2_ifu_mem_ctl.scala 426:70]
  wire  _T_1508 = _T_1506 & _T_58; // @[el2_ifu_mem_ctl.scala 426:92]
  wire  _T_1509 = _T_1502 | _T_1508; // @[el2_ifu_mem_ctl.scala 425:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 428:58]
  wire  _T_1510 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 427:28]
  wire  _T_1511 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 427:50]
  wire  _T_1512 = _T_1510 & _T_1511; // @[el2_ifu_mem_ctl.scala 427:48]
  wire  _T_1514 = _T_1512 & _T_319; // @[el2_ifu_mem_ctl.scala 427:70]
  wire  ic_crit_wd_rdy_new_in = _T_1509 | _T_1514; // @[el2_ifu_mem_ctl.scala 426:117]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 629:43]
  wire  _T_1251 = ic_crit_wd_rdy | _T_2219; // @[el2_ifu_mem_ctl.scala 372:38]
  wire  _T_1253 = _T_1251 | _T_2235; // @[el2_ifu_mem_ctl.scala 372:64]
  wire  _T_1254 = ~_T_1253; // @[el2_ifu_mem_ctl.scala 372:21]
  wire  _T_1255 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 372:98]
  wire  sel_ic_data = _T_1254 & _T_1255; // @[el2_ifu_mem_ctl.scala 372:96]
  wire  _T_2442 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 472:44]
  wire  _T_1608 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 439:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 411:60]
  wire  _T_1552 = _T_1399 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1553 = _T_1402 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1560 = _T_1552 | _T_1553; // @[Mux.scala 27:72]
  wire  _T_1554 = _T_1405 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1561 = _T_1560 | _T_1554; // @[Mux.scala 27:72]
  wire  _T_1555 = _T_1408 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1562 = _T_1561 | _T_1555; // @[Mux.scala 27:72]
  wire  _T_1556 = _T_1411 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1563 = _T_1562 | _T_1556; // @[Mux.scala 27:72]
  wire  _T_1557 = _T_1414 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1564 = _T_1563 | _T_1557; // @[Mux.scala 27:72]
  wire  _T_1558 = _T_1417 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1565 = _T_1564 | _T_1558; // @[Mux.scala 27:72]
  wire  _T_1559 = _T_1420 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1565 | _T_1559; // @[Mux.scala 27:72]
  wire  _T_1591 = _T_2152 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1592 = _T_2155 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1599 = _T_1591 | _T_1592; // @[Mux.scala 27:72]
  wire  _T_1593 = _T_2158 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1600 = _T_1599 | _T_1593; // @[Mux.scala 27:72]
  wire  _T_1594 = _T_2161 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1601 = _T_1600 | _T_1594; // @[Mux.scala 27:72]
  wire  _T_1595 = _T_2164 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1602 = _T_1601 | _T_1595; // @[Mux.scala 27:72]
  wire  _T_1596 = _T_2167 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1603 = _T_1602 | _T_1596; // @[Mux.scala 27:72]
  wire  _T_1597 = _T_2170 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1604 = _T_1603 | _T_1597; // @[Mux.scala 27:72]
  wire  _T_1598 = _T_2173 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1604 | _T_1598; // @[Mux.scala 27:72]
  wire  _T_1609 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 441:70]
  wire  ifu_byp_data_err_new = _T_1608 ? ic_miss_buff_data_error_bypass : _T_1609; // @[el2_ifu_mem_ctl.scala 439:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 383:42]
  wire  _T_2443 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 472:91]
  wire  _T_2444 = ~_T_2443; // @[el2_ifu_mem_ctl.scala 472:60]
  wire  ic_rd_parity_final_err = _T_2442 & _T_2444; // @[el2_ifu_mem_ctl.scala 472:58]
  reg  ic_debug_ict_array_sel_ff; // @[el2_ifu_mem_ctl.scala 837:63]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9323 = _T_4620 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 764:8]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9325 = _T_4621 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9578 = _T_9323 | _T_9325; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9327 = _T_4622 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9579 = _T_9578 | _T_9327; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9329 = _T_4623 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9580 = _T_9579 | _T_9329; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9331 = _T_4624 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9581 = _T_9580 | _T_9331; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9333 = _T_4625 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9582 = _T_9581 | _T_9333; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9335 = _T_4626 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9583 = _T_9582 | _T_9335; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9337 = _T_4627 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9584 = _T_9583 | _T_9337; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9339 = _T_4628 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9585 = _T_9584 | _T_9339; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9341 = _T_4629 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9586 = _T_9585 | _T_9341; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9343 = _T_4630 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9587 = _T_9586 | _T_9343; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9345 = _T_4631 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9588 = _T_9587 | _T_9345; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9347 = _T_4632 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9589 = _T_9588 | _T_9347; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9349 = _T_4633 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9590 = _T_9589 | _T_9349; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9351 = _T_4634 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9591 = _T_9590 | _T_9351; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9353 = _T_4635 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9592 = _T_9591 | _T_9353; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9355 = _T_4636 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9593 = _T_9592 | _T_9355; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9357 = _T_4637 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9594 = _T_9593 | _T_9357; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9359 = _T_4638 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9595 = _T_9594 | _T_9359; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9361 = _T_4639 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9596 = _T_9595 | _T_9361; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9363 = _T_4640 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9597 = _T_9596 | _T_9363; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9365 = _T_4641 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9598 = _T_9597 | _T_9365; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9367 = _T_4642 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9599 = _T_9598 | _T_9367; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9369 = _T_4643 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9600 = _T_9599 | _T_9369; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9371 = _T_4644 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9601 = _T_9600 | _T_9371; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9373 = _T_4645 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9602 = _T_9601 | _T_9373; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9375 = _T_4646 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9603 = _T_9602 | _T_9375; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9377 = _T_4647 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9604 = _T_9603 | _T_9377; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9379 = _T_4648 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9605 = _T_9604 | _T_9379; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9381 = _T_4649 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9606 = _T_9605 | _T_9381; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9383 = _T_4650 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9607 = _T_9606 | _T_9383; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9385 = _T_4651 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9608 = _T_9607 | _T_9385; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9387 = _T_4652 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9609 = _T_9608 | _T_9387; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9389 = _T_4653 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9610 = _T_9609 | _T_9389; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9391 = _T_4654 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9611 = _T_9610 | _T_9391; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9393 = _T_4655 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9612 = _T_9611 | _T_9393; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9395 = _T_4656 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9613 = _T_9612 | _T_9395; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9397 = _T_4657 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9614 = _T_9613 | _T_9397; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9399 = _T_4658 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9615 = _T_9614 | _T_9399; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9401 = _T_4659 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9616 = _T_9615 | _T_9401; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9403 = _T_4660 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9617 = _T_9616 | _T_9403; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9405 = _T_4661 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9618 = _T_9617 | _T_9405; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9407 = _T_4662 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9619 = _T_9618 | _T_9407; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9409 = _T_4663 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9620 = _T_9619 | _T_9409; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9411 = _T_4664 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9621 = _T_9620 | _T_9411; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9413 = _T_4665 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9622 = _T_9621 | _T_9413; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9415 = _T_4666 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9623 = _T_9622 | _T_9415; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9417 = _T_4667 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9624 = _T_9623 | _T_9417; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9419 = _T_4668 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9625 = _T_9624 | _T_9419; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9421 = _T_4669 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9626 = _T_9625 | _T_9421; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9423 = _T_4670 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9627 = _T_9626 | _T_9423; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9425 = _T_4671 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9628 = _T_9627 | _T_9425; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9427 = _T_4672 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9629 = _T_9628 | _T_9427; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9429 = _T_4673 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9630 = _T_9629 | _T_9429; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9431 = _T_4674 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9631 = _T_9630 | _T_9431; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9433 = _T_4675 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9632 = _T_9631 | _T_9433; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9435 = _T_4676 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9633 = _T_9632 | _T_9435; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9437 = _T_4677 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9634 = _T_9633 | _T_9437; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9439 = _T_4678 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9635 = _T_9634 | _T_9439; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9441 = _T_4679 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9636 = _T_9635 | _T_9441; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9443 = _T_4680 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9637 = _T_9636 | _T_9443; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9445 = _T_4681 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9638 = _T_9637 | _T_9445; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9447 = _T_4682 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9639 = _T_9638 | _T_9447; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9449 = _T_4683 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9640 = _T_9639 | _T_9449; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9451 = _T_4684 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9641 = _T_9640 | _T_9451; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9453 = _T_4685 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9642 = _T_9641 | _T_9453; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9455 = _T_4686 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9643 = _T_9642 | _T_9455; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9457 = _T_4687 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9644 = _T_9643 | _T_9457; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9459 = _T_4688 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9645 = _T_9644 | _T_9459; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9461 = _T_4689 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9646 = _T_9645 | _T_9461; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9463 = _T_4690 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9647 = _T_9646 | _T_9463; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9465 = _T_4691 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9648 = _T_9647 | _T_9465; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9467 = _T_4692 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9649 = _T_9648 | _T_9467; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9469 = _T_4693 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9650 = _T_9649 | _T_9469; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9471 = _T_4694 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9651 = _T_9650 | _T_9471; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9473 = _T_4695 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9652 = _T_9651 | _T_9473; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9475 = _T_4696 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9653 = _T_9652 | _T_9475; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9477 = _T_4697 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9654 = _T_9653 | _T_9477; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9479 = _T_4698 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9655 = _T_9654 | _T_9479; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9481 = _T_4699 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9656 = _T_9655 | _T_9481; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9483 = _T_4700 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9657 = _T_9656 | _T_9483; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9485 = _T_4701 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9658 = _T_9657 | _T_9485; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9487 = _T_4702 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9659 = _T_9658 | _T_9487; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9489 = _T_4703 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9660 = _T_9659 | _T_9489; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9491 = _T_4704 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9661 = _T_9660 | _T_9491; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9493 = _T_4705 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9662 = _T_9661 | _T_9493; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9495 = _T_4706 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9663 = _T_9662 | _T_9495; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9497 = _T_4707 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9664 = _T_9663 | _T_9497; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9499 = _T_4708 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9665 = _T_9664 | _T_9499; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9501 = _T_4709 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9666 = _T_9665 | _T_9501; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9503 = _T_4710 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9667 = _T_9666 | _T_9503; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9505 = _T_4711 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9668 = _T_9667 | _T_9505; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9507 = _T_4712 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9669 = _T_9668 | _T_9507; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9509 = _T_4713 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9670 = _T_9669 | _T_9509; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9511 = _T_4714 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9671 = _T_9670 | _T_9511; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9513 = _T_4715 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9672 = _T_9671 | _T_9513; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9515 = _T_4716 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9673 = _T_9672 | _T_9515; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9517 = _T_4717 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9674 = _T_9673 | _T_9517; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9519 = _T_4718 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9675 = _T_9674 | _T_9519; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9521 = _T_4719 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9676 = _T_9675 | _T_9521; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9523 = _T_4720 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9677 = _T_9676 | _T_9523; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9525 = _T_4721 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9678 = _T_9677 | _T_9525; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9527 = _T_4722 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9679 = _T_9678 | _T_9527; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9529 = _T_4723 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9680 = _T_9679 | _T_9529; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9531 = _T_4724 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9681 = _T_9680 | _T_9531; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9533 = _T_4725 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9682 = _T_9681 | _T_9533; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9535 = _T_4726 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9683 = _T_9682 | _T_9535; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9537 = _T_4727 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9684 = _T_9683 | _T_9537; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9539 = _T_4728 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9685 = _T_9684 | _T_9539; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9541 = _T_4729 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9686 = _T_9685 | _T_9541; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9543 = _T_4730 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9687 = _T_9686 | _T_9543; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9545 = _T_4731 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9688 = _T_9687 | _T_9545; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9547 = _T_4732 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9689 = _T_9688 | _T_9547; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9549 = _T_4733 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9690 = _T_9689 | _T_9549; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9551 = _T_4734 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9691 = _T_9690 | _T_9551; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9553 = _T_4735 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9692 = _T_9691 | _T_9553; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9555 = _T_4736 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9693 = _T_9692 | _T_9555; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9557 = _T_4737 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9694 = _T_9693 | _T_9557; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9559 = _T_4738 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9695 = _T_9694 | _T_9559; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9561 = _T_4739 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9696 = _T_9695 | _T_9561; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9563 = _T_4740 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9697 = _T_9696 | _T_9563; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9565 = _T_4741 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9698 = _T_9697 | _T_9565; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9567 = _T_4742 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9699 = _T_9698 | _T_9567; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9569 = _T_4743 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9700 = _T_9699 | _T_9569; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9571 = _T_4744 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9701 = _T_9700 | _T_9571; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9573 = _T_4745 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9702 = _T_9701 | _T_9573; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9575 = _T_4746 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9703 = _T_9702 | _T_9575; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9577 = _T_4747 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9704 = _T_9703 | _T_9577; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8940 = _T_4620 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 764:8]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8942 = _T_4621 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9195 = _T_8940 | _T_8942; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8944 = _T_4622 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9196 = _T_9195 | _T_8944; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8946 = _T_4623 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9197 = _T_9196 | _T_8946; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8948 = _T_4624 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9198 = _T_9197 | _T_8948; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_8950 = _T_4625 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9199 = _T_9198 | _T_8950; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_8952 = _T_4626 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9200 = _T_9199 | _T_8952; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_8954 = _T_4627 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9201 = _T_9200 | _T_8954; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_8956 = _T_4628 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9202 = _T_9201 | _T_8956; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_8958 = _T_4629 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9203 = _T_9202 | _T_8958; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_8960 = _T_4630 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9204 = _T_9203 | _T_8960; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_8962 = _T_4631 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9205 = _T_9204 | _T_8962; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_8964 = _T_4632 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9206 = _T_9205 | _T_8964; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_8966 = _T_4633 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9207 = _T_9206 | _T_8966; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_8968 = _T_4634 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9208 = _T_9207 | _T_8968; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_8970 = _T_4635 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9209 = _T_9208 | _T_8970; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_8972 = _T_4636 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9210 = _T_9209 | _T_8972; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_8974 = _T_4637 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9211 = _T_9210 | _T_8974; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_8976 = _T_4638 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9212 = _T_9211 | _T_8976; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_8978 = _T_4639 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9213 = _T_9212 | _T_8978; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_8980 = _T_4640 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9214 = _T_9213 | _T_8980; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_8982 = _T_4641 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9215 = _T_9214 | _T_8982; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_8984 = _T_4642 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9216 = _T_9215 | _T_8984; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_8986 = _T_4643 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9217 = _T_9216 | _T_8986; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_8988 = _T_4644 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9218 = _T_9217 | _T_8988; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_8990 = _T_4645 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9219 = _T_9218 | _T_8990; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_8992 = _T_4646 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9220 = _T_9219 | _T_8992; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_8994 = _T_4647 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9221 = _T_9220 | _T_8994; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_8996 = _T_4648 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9222 = _T_9221 | _T_8996; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_8998 = _T_4649 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9223 = _T_9222 | _T_8998; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9000 = _T_4650 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9224 = _T_9223 | _T_9000; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9002 = _T_4651 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9225 = _T_9224 | _T_9002; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9004 = _T_4652 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9226 = _T_9225 | _T_9004; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9006 = _T_4653 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9227 = _T_9226 | _T_9006; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9008 = _T_4654 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9228 = _T_9227 | _T_9008; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9010 = _T_4655 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9229 = _T_9228 | _T_9010; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9012 = _T_4656 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9230 = _T_9229 | _T_9012; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9014 = _T_4657 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9231 = _T_9230 | _T_9014; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9016 = _T_4658 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9232 = _T_9231 | _T_9016; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9018 = _T_4659 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9233 = _T_9232 | _T_9018; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9020 = _T_4660 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9234 = _T_9233 | _T_9020; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9022 = _T_4661 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9235 = _T_9234 | _T_9022; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9024 = _T_4662 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9236 = _T_9235 | _T_9024; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9026 = _T_4663 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9237 = _T_9236 | _T_9026; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9028 = _T_4664 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9238 = _T_9237 | _T_9028; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9030 = _T_4665 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9239 = _T_9238 | _T_9030; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9032 = _T_4666 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9240 = _T_9239 | _T_9032; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9034 = _T_4667 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9241 = _T_9240 | _T_9034; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9036 = _T_4668 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9242 = _T_9241 | _T_9036; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9038 = _T_4669 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9243 = _T_9242 | _T_9038; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9040 = _T_4670 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9244 = _T_9243 | _T_9040; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9042 = _T_4671 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9245 = _T_9244 | _T_9042; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9044 = _T_4672 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9246 = _T_9245 | _T_9044; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9046 = _T_4673 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9247 = _T_9246 | _T_9046; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9048 = _T_4674 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9248 = _T_9247 | _T_9048; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9050 = _T_4675 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9249 = _T_9248 | _T_9050; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9052 = _T_4676 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9250 = _T_9249 | _T_9052; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9054 = _T_4677 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9251 = _T_9250 | _T_9054; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9056 = _T_4678 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9252 = _T_9251 | _T_9056; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9058 = _T_4679 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9253 = _T_9252 | _T_9058; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9060 = _T_4680 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9254 = _T_9253 | _T_9060; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9062 = _T_4681 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9255 = _T_9254 | _T_9062; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9064 = _T_4682 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9256 = _T_9255 | _T_9064; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9066 = _T_4683 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9257 = _T_9256 | _T_9066; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9068 = _T_4684 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9258 = _T_9257 | _T_9068; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9070 = _T_4685 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9259 = _T_9258 | _T_9070; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9072 = _T_4686 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9260 = _T_9259 | _T_9072; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9074 = _T_4687 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9261 = _T_9260 | _T_9074; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9076 = _T_4688 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9262 = _T_9261 | _T_9076; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9078 = _T_4689 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9263 = _T_9262 | _T_9078; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9080 = _T_4690 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9264 = _T_9263 | _T_9080; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9082 = _T_4691 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9265 = _T_9264 | _T_9082; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9084 = _T_4692 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9266 = _T_9265 | _T_9084; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9086 = _T_4693 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9267 = _T_9266 | _T_9086; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9088 = _T_4694 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9268 = _T_9267 | _T_9088; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9090 = _T_4695 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9269 = _T_9268 | _T_9090; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9092 = _T_4696 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9270 = _T_9269 | _T_9092; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9094 = _T_4697 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9271 = _T_9270 | _T_9094; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9096 = _T_4698 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9272 = _T_9271 | _T_9096; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9098 = _T_4699 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9273 = _T_9272 | _T_9098; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9100 = _T_4700 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9274 = _T_9273 | _T_9100; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9102 = _T_4701 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9275 = _T_9274 | _T_9102; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9104 = _T_4702 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9276 = _T_9275 | _T_9104; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9106 = _T_4703 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9277 = _T_9276 | _T_9106; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9108 = _T_4704 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9278 = _T_9277 | _T_9108; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9110 = _T_4705 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9279 = _T_9278 | _T_9110; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9112 = _T_4706 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9280 = _T_9279 | _T_9112; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9114 = _T_4707 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9281 = _T_9280 | _T_9114; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9116 = _T_4708 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9282 = _T_9281 | _T_9116; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9118 = _T_4709 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9283 = _T_9282 | _T_9118; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9120 = _T_4710 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9284 = _T_9283 | _T_9120; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9122 = _T_4711 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9285 = _T_9284 | _T_9122; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9124 = _T_4712 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9286 = _T_9285 | _T_9124; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9126 = _T_4713 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9287 = _T_9286 | _T_9126; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9128 = _T_4714 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9288 = _T_9287 | _T_9128; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9130 = _T_4715 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9289 = _T_9288 | _T_9130; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9132 = _T_4716 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9290 = _T_9289 | _T_9132; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9134 = _T_4717 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9291 = _T_9290 | _T_9134; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9136 = _T_4718 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9292 = _T_9291 | _T_9136; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9138 = _T_4719 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9293 = _T_9292 | _T_9138; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9140 = _T_4720 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9294 = _T_9293 | _T_9140; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9142 = _T_4721 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9295 = _T_9294 | _T_9142; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9144 = _T_4722 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9296 = _T_9295 | _T_9144; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9146 = _T_4723 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9297 = _T_9296 | _T_9146; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9148 = _T_4724 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9298 = _T_9297 | _T_9148; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9150 = _T_4725 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9299 = _T_9298 | _T_9150; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9152 = _T_4726 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9300 = _T_9299 | _T_9152; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9154 = _T_4727 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9301 = _T_9300 | _T_9154; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9156 = _T_4728 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9302 = _T_9301 | _T_9156; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9158 = _T_4729 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9303 = _T_9302 | _T_9158; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9160 = _T_4730 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9304 = _T_9303 | _T_9160; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9162 = _T_4731 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9305 = _T_9304 | _T_9162; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9164 = _T_4732 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9306 = _T_9305 | _T_9164; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9166 = _T_4733 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9307 = _T_9306 | _T_9166; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9168 = _T_4734 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9308 = _T_9307 | _T_9168; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9170 = _T_4735 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9309 = _T_9308 | _T_9170; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9172 = _T_4736 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9310 = _T_9309 | _T_9172; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9174 = _T_4737 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9311 = _T_9310 | _T_9174; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9176 = _T_4738 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9312 = _T_9311 | _T_9176; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9178 = _T_4739 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9313 = _T_9312 | _T_9178; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9180 = _T_4740 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9314 = _T_9313 | _T_9180; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9182 = _T_4741 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9315 = _T_9314 | _T_9182; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9184 = _T_4742 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9316 = _T_9315 | _T_9184; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9186 = _T_4743 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9317 = _T_9316 | _T_9186; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9188 = _T_4744 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9318 = _T_9317 | _T_9188; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9190 = _T_4745 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9319 = _T_9318 | _T_9190; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9192 = _T_4746 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9320 = _T_9319 | _T_9192; // @[el2_ifu_mem_ctl.scala 764:89]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9194 = _T_4747 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 764:8]
  wire  _T_9321 = _T_9320 | _T_9194; // @[el2_ifu_mem_ctl.scala 764:89]
  wire [1:0] ic_tag_valid_unq = {_T_9704,_T_9321}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[el2_ifu_mem_ctl.scala 836:53]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 838:54]
  wire [1:0] _T_9744 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9745 = ic_debug_way_ff & _T_9744; // @[el2_ifu_mem_ctl.scala 819:67]
  wire [1:0] _T_9746 = ic_tag_valid_unq & _T_9745; // @[el2_ifu_mem_ctl.scala 819:48]
  wire  ic_debug_tag_val_rd_out = |_T_9746; // @[el2_ifu_mem_ctl.scala 819:115]
  wire [70:0] _T_1210 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],6'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1211; // @[el2_ifu_mem_ctl.scala 355:63]
  wire  _T_1249 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 371:98]
  wire  sel_byp_data = _T_1253 & _T_1249; // @[el2_ifu_mem_ctl.scala 371:96]
  wire [63:0] _T_1260 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1261 = _T_1260 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 378:69]
  wire [63:0] _T_1263 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2099 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 447:31]
  wire  _T_1612 = ~ifu_fetch_addr_int_f[1]; // @[el2_ifu_mem_ctl.scala 443:38]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1613 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1661 = _T_1613 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1616 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1662 = _T_1616 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1677 = _T_1661 | _T_1662; // @[Mux.scala 27:72]
  wire  _T_1619 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1663 = _T_1619 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1678 = _T_1677 | _T_1663; // @[Mux.scala 27:72]
  wire  _T_1622 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1664 = _T_1622 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1679 = _T_1678 | _T_1664; // @[Mux.scala 27:72]
  wire  _T_1625 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1665 = _T_1625 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1680 = _T_1679 | _T_1665; // @[Mux.scala 27:72]
  wire  _T_1628 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1666 = _T_1628 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1681 = _T_1680 | _T_1666; // @[Mux.scala 27:72]
  wire  _T_1631 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1667 = _T_1631 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1682 = _T_1681 | _T_1667; // @[Mux.scala 27:72]
  wire  _T_1634 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1668 = _T_1634 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1683 = _T_1682 | _T_1668; // @[Mux.scala 27:72]
  wire  _T_1637 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1669 = _T_1637 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1684 = _T_1683 | _T_1669; // @[Mux.scala 27:72]
  wire  _T_1640 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1670 = _T_1640 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1685 = _T_1684 | _T_1670; // @[Mux.scala 27:72]
  wire  _T_1643 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1671 = _T_1643 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1686 = _T_1685 | _T_1671; // @[Mux.scala 27:72]
  wire  _T_1646 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1672 = _T_1646 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1687 = _T_1686 | _T_1672; // @[Mux.scala 27:72]
  wire  _T_1649 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1673 = _T_1649 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1688 = _T_1687 | _T_1673; // @[Mux.scala 27:72]
  wire  _T_1652 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1674 = _T_1652 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1689 = _T_1688 | _T_1674; // @[Mux.scala 27:72]
  wire  _T_1655 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1675 = _T_1655 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1690 = _T_1689 | _T_1675; // @[Mux.scala 27:72]
  wire  _T_1658 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 444:73]
  wire [15:0] _T_1676 = _T_1658 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1691 = _T_1690 | _T_1676; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1693 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1741 = _T_1693 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1696 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1742 = _T_1696 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1757 = _T_1741 | _T_1742; // @[Mux.scala 27:72]
  wire  _T_1699 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1743 = _T_1699 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1758 = _T_1757 | _T_1743; // @[Mux.scala 27:72]
  wire  _T_1702 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1744 = _T_1702 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1759 = _T_1758 | _T_1744; // @[Mux.scala 27:72]
  wire  _T_1705 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1745 = _T_1705 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1760 = _T_1759 | _T_1745; // @[Mux.scala 27:72]
  wire  _T_1708 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1746 = _T_1708 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1761 = _T_1760 | _T_1746; // @[Mux.scala 27:72]
  wire  _T_1711 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1747 = _T_1711 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1762 = _T_1761 | _T_1747; // @[Mux.scala 27:72]
  wire  _T_1714 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1748 = _T_1714 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1763 = _T_1762 | _T_1748; // @[Mux.scala 27:72]
  wire  _T_1717 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1749 = _T_1717 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1764 = _T_1763 | _T_1749; // @[Mux.scala 27:72]
  wire  _T_1720 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1750 = _T_1720 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1765 = _T_1764 | _T_1750; // @[Mux.scala 27:72]
  wire  _T_1723 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1751 = _T_1723 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1766 = _T_1765 | _T_1751; // @[Mux.scala 27:72]
  wire  _T_1726 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1752 = _T_1726 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1767 = _T_1766 | _T_1752; // @[Mux.scala 27:72]
  wire  _T_1729 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1753 = _T_1729 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1768 = _T_1767 | _T_1753; // @[Mux.scala 27:72]
  wire  _T_1732 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1754 = _T_1732 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1769 = _T_1768 | _T_1754; // @[Mux.scala 27:72]
  wire  _T_1735 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1755 = _T_1735 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1770 = _T_1769 | _T_1755; // @[Mux.scala 27:72]
  wire  _T_1738 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 444:179]
  wire [31:0] _T_1756 = _T_1738 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1771 = _T_1770 | _T_1756; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1773 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1821 = _T_1773 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1776 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1822 = _T_1776 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1837 = _T_1821 | _T_1822; // @[Mux.scala 27:72]
  wire  _T_1779 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1823 = _T_1779 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1838 = _T_1837 | _T_1823; // @[Mux.scala 27:72]
  wire  _T_1782 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1824 = _T_1782 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1839 = _T_1838 | _T_1824; // @[Mux.scala 27:72]
  wire  _T_1785 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1825 = _T_1785 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1840 = _T_1839 | _T_1825; // @[Mux.scala 27:72]
  wire  _T_1788 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1826 = _T_1788 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1841 = _T_1840 | _T_1826; // @[Mux.scala 27:72]
  wire  _T_1791 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1827 = _T_1791 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1842 = _T_1841 | _T_1827; // @[Mux.scala 27:72]
  wire  _T_1794 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1828 = _T_1794 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1843 = _T_1842 | _T_1828; // @[Mux.scala 27:72]
  wire  _T_1797 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1829 = _T_1797 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1844 = _T_1843 | _T_1829; // @[Mux.scala 27:72]
  wire  _T_1800 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1830 = _T_1800 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1845 = _T_1844 | _T_1830; // @[Mux.scala 27:72]
  wire  _T_1803 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1831 = _T_1803 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1846 = _T_1845 | _T_1831; // @[Mux.scala 27:72]
  wire  _T_1806 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1832 = _T_1806 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1847 = _T_1846 | _T_1832; // @[Mux.scala 27:72]
  wire  _T_1809 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1833 = _T_1809 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1848 = _T_1847 | _T_1833; // @[Mux.scala 27:72]
  wire  _T_1812 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1834 = _T_1812 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1849 = _T_1848 | _T_1834; // @[Mux.scala 27:72]
  wire  _T_1815 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1835 = _T_1815 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1850 = _T_1849 | _T_1835; // @[Mux.scala 27:72]
  wire  _T_1818 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 444:285]
  wire [31:0] _T_1836 = _T_1818 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1851 = _T_1850 | _T_1836; // @[Mux.scala 27:72]
  wire [79:0] _T_1854 = {_T_1691,_T_1771,_T_1851}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1855 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1903 = _T_1855 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1858 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1904 = _T_1858 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1919 = _T_1903 | _T_1904; // @[Mux.scala 27:72]
  wire  _T_1861 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1905 = _T_1861 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1920 = _T_1919 | _T_1905; // @[Mux.scala 27:72]
  wire  _T_1864 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1906 = _T_1864 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1921 = _T_1920 | _T_1906; // @[Mux.scala 27:72]
  wire  _T_1867 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1907 = _T_1867 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1922 = _T_1921 | _T_1907; // @[Mux.scala 27:72]
  wire  _T_1870 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1908 = _T_1870 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1923 = _T_1922 | _T_1908; // @[Mux.scala 27:72]
  wire  _T_1873 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1909 = _T_1873 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1924 = _T_1923 | _T_1909; // @[Mux.scala 27:72]
  wire  _T_1876 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1910 = _T_1876 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1925 = _T_1924 | _T_1910; // @[Mux.scala 27:72]
  wire  _T_1879 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1911 = _T_1879 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1926 = _T_1925 | _T_1911; // @[Mux.scala 27:72]
  wire  _T_1882 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1912 = _T_1882 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1927 = _T_1926 | _T_1912; // @[Mux.scala 27:72]
  wire  _T_1885 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1913 = _T_1885 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1928 = _T_1927 | _T_1913; // @[Mux.scala 27:72]
  wire  _T_1888 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1914 = _T_1888 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1929 = _T_1928 | _T_1914; // @[Mux.scala 27:72]
  wire  _T_1891 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1915 = _T_1891 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1930 = _T_1929 | _T_1915; // @[Mux.scala 27:72]
  wire  _T_1894 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1916 = _T_1894 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1931 = _T_1930 | _T_1916; // @[Mux.scala 27:72]
  wire  _T_1897 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1917 = _T_1897 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1932 = _T_1931 | _T_1917; // @[Mux.scala 27:72]
  wire  _T_1900 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1918 = _T_1900 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1933 = _T_1932 | _T_1918; // @[Mux.scala 27:72]
  wire [31:0] _T_1983 = _T_1613 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1984 = _T_1616 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1983 | _T_1984; // @[Mux.scala 27:72]
  wire [31:0] _T_1985 = _T_1619 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1999 | _T_1985; // @[Mux.scala 27:72]
  wire [31:0] _T_1986 = _T_1622 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_2000 | _T_1986; // @[Mux.scala 27:72]
  wire [31:0] _T_1987 = _T_1625 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_2001 | _T_1987; // @[Mux.scala 27:72]
  wire [31:0] _T_1988 = _T_1628 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_2002 | _T_1988; // @[Mux.scala 27:72]
  wire [31:0] _T_1989 = _T_1631 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_2003 | _T_1989; // @[Mux.scala 27:72]
  wire [31:0] _T_1990 = _T_1634 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_2004 | _T_1990; // @[Mux.scala 27:72]
  wire [31:0] _T_1991 = _T_1637 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_2005 | _T_1991; // @[Mux.scala 27:72]
  wire [31:0] _T_1992 = _T_1640 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_2006 | _T_1992; // @[Mux.scala 27:72]
  wire [31:0] _T_1993 = _T_1643 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_2007 | _T_1993; // @[Mux.scala 27:72]
  wire [31:0] _T_1994 = _T_1646 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_2008 | _T_1994; // @[Mux.scala 27:72]
  wire [31:0] _T_1995 = _T_1649 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_2009 | _T_1995; // @[Mux.scala 27:72]
  wire [31:0] _T_1996 = _T_1652 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_2010 | _T_1996; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1655 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_2011 | _T_1997; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1658 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_2012 | _T_1998; // @[Mux.scala 27:72]
  wire [79:0] _T_2096 = {_T_1933,_T_2013,_T_1771}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1612 ? _T_1854 : _T_2096; // @[el2_ifu_mem_ctl.scala 443:37]
  wire [79:0] _T_2101 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2099 ? ic_byp_data_only_pre_new : _T_2101; // @[el2_ifu_mem_ctl.scala 447:30]
  wire [79:0] _GEN_447 = {{16'd0}, _T_1263}; // @[el2_ifu_mem_ctl.scala 378:114]
  wire [79:0] _T_1264 = _GEN_447 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 378:114]
  wire [79:0] _GEN_448 = {{16'd0}, _T_1261}; // @[el2_ifu_mem_ctl.scala 378:88]
  wire [79:0] ic_premux_data_temp = _GEN_448 | _T_1264; // @[el2_ifu_mem_ctl.scala 378:88]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_319; // @[el2_ifu_mem_ctl.scala 385:38]
  reg  ifc_region_acc_fault_memory_f; // @[el2_ifu_mem_ctl.scala 851:66]
  wire [1:0] _T_1272 = ifc_region_acc_fault_memory_f ? 2'h3 : 2'h0; // @[el2_ifu_mem_ctl.scala 390:10]
  wire [1:0] _T_1273 = ifc_region_acc_fault_f ? 2'h2 : _T_1272; // @[el2_ifu_mem_ctl.scala 389:8]
  wire  _T_1275 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[el2_ifu_mem_ctl.scala 391:45]
  wire  _T_1277 = byp_fetch_index == 5'h1f; // @[el2_ifu_mem_ctl.scala 391:80]
  wire  _T_1278 = ~_T_1277; // @[el2_ifu_mem_ctl.scala 391:71]
  wire  _T_1279 = _T_1275 & _T_1278; // @[el2_ifu_mem_ctl.scala 391:69]
  wire  _T_1280 = err_stop_state != 2'h2; // @[el2_ifu_mem_ctl.scala 391:131]
  wire  _T_1281 = _T_1279 & _T_1280; // @[el2_ifu_mem_ctl.scala 391:114]
  wire [6:0] _T_1353 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1}; // @[Cat.scala 29:58]
  wire  _T_1359 = ic_miss_buff_data_error[0] & _T_1325; // @[el2_ifu_mem_ctl.scala 410:32]
  wire  _T_2641 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 625:47]
  wire  _T_2642 = _T_2641 & _T_13; // @[el2_ifu_mem_ctl.scala 625:50]
  wire  bus_ifu_wr_data_error = _T_2642 & miss_pending; // @[el2_ifu_mem_ctl.scala 625:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1359; // @[el2_ifu_mem_ctl.scala 409:72]
  wire  _T_1363 = ic_miss_buff_data_error[1] & _T_1325; // @[el2_ifu_mem_ctl.scala 410:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1363; // @[el2_ifu_mem_ctl.scala 409:72]
  wire  _T_1367 = ic_miss_buff_data_error[2] & _T_1325; // @[el2_ifu_mem_ctl.scala 410:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1367; // @[el2_ifu_mem_ctl.scala 409:72]
  wire  _T_1371 = ic_miss_buff_data_error[3] & _T_1325; // @[el2_ifu_mem_ctl.scala 410:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1371; // @[el2_ifu_mem_ctl.scala 409:72]
  wire  _T_1375 = ic_miss_buff_data_error[4] & _T_1325; // @[el2_ifu_mem_ctl.scala 410:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1375; // @[el2_ifu_mem_ctl.scala 409:72]
  wire  _T_1379 = ic_miss_buff_data_error[5] & _T_1325; // @[el2_ifu_mem_ctl.scala 410:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1379; // @[el2_ifu_mem_ctl.scala 409:72]
  wire  _T_1383 = ic_miss_buff_data_error[6] & _T_1325; // @[el2_ifu_mem_ctl.scala 410:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1383; // @[el2_ifu_mem_ctl.scala 409:72]
  wire  _T_1387 = ic_miss_buff_data_error[7] & _T_1325; // @[el2_ifu_mem_ctl.scala 410:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1387; // @[el2_ifu_mem_ctl.scala 409:72]
  wire [6:0] _T_1393 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1}; // @[Cat.scala 29:58]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2451 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2459 = _T_6 & _T_319; // @[el2_ifu_mem_ctl.scala 492:65]
  wire  _T_2460 = _T_2459 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 492:88]
  wire  _T_2462 = _T_2460 & _T_2574; // @[el2_ifu_mem_ctl.scala 492:112]
  wire  _T_2463 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2464 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 497:50]
  wire  _T_2466 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2473 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2475 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_22 = _T_2473 | _T_2475; // @[Conditional.scala 39:67]
  wire  _GEN_24 = _T_2466 ? _T_2464 : _GEN_22; // @[Conditional.scala 39:67]
  wire  _GEN_26 = _T_2463 ? _T_2464 : _GEN_24; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2451 ? _T_2462 : _GEN_26; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2451 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2465 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 498:56]
  wire  _GEN_27 = _T_2463 & _T_2465; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2451 ? 1'h0 : _GEN_27; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 483:58]
  wire  _T_2448 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 482:49]
  wire  _T_2453 = io_ic_error_start & _T_319; // @[el2_ifu_mem_ctl.scala 491:87]
  wire  _T_2467 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 501:30]
  wire  _T_2468 = _T_2467 & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 501:55]
  wire  _T_2469 = _T_2468 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 501:85]
  wire  _T_2478 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 522:66]
  wire  _T_2479 = io_dec_tlu_flush_err_wb & _T_2478; // @[el2_ifu_mem_ctl.scala 522:52]
  wire  _T_2481 = _T_2479 & _T_2574; // @[el2_ifu_mem_ctl.scala 522:81]
  wire  _T_2483 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 525:59]
  wire  _T_2484 = _T_2483 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 525:86]
  wire  _T_2498 = _T_2483 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 528:81]
  wire  _T_2499 = _T_2498 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 528:103]
  wire  _T_2500 = _T_2499 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 528:126]
  wire  _T_2520 = _T_2498 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 535:103]
  wire  _T_2528 = io_dec_tlu_flush_lower_wb & _T_2467; // @[el2_ifu_mem_ctl.scala 540:60]
  wire  _T_2529 = _T_2528 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 540:88]
  wire  _T_2530 = _T_2529 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 540:115]
  wire  _GEN_34 = _T_2526 & _T_2484; // @[Conditional.scala 39:67]
  wire  _GEN_37 = _T_2509 ? _T_2520 : _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_39 = _T_2509 | _T_2526; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_2482 ? _T_2500 : _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_2482 | _GEN_39; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2477 ? _T_2481 : _GEN_41; // @[Conditional.scala 40:58]
  reg  bus_cmd_req_hold; // @[el2_ifu_mem_ctl.scala 563:53]
  wire  _T_2542 = ic_act_miss_f | bus_cmd_req_hold; // @[el2_ifu_mem_ctl.scala 559:45]
  reg  ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 560:55]
  wire  _T_2543 = _T_2542 | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 559:64]
  wire  _T_2545 = _T_2543 & _T_2574; // @[el2_ifu_mem_ctl.scala 559:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2547 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 559:133]
  wire  _T_2548 = _T_2547 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 559:164]
  wire  _T_2549 = _T_2548 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 559:184]
  wire  _T_2550 = _T_2549 & miss_pending; // @[el2_ifu_mem_ctl.scala 559:204]
  wire  _T_2551 = ~_T_2550; // @[el2_ifu_mem_ctl.scala 559:112]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 591:45]
  wire  _T_2568 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 594:35]
  wire  _T_2569 = _T_2568 & miss_pending; // @[el2_ifu_mem_ctl.scala 594:53]
  wire  bus_cmd_sent = _T_2569 & _T_2574; // @[el2_ifu_mem_ctl.scala 594:68]
  wire  _T_2554 = ~bus_cmd_sent; // @[el2_ifu_mem_ctl.scala 562:61]
  wire  _T_2555 = _T_2542 & _T_2554; // @[el2_ifu_mem_ctl.scala 562:59]
  wire [2:0] _T_2559 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2561 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2563 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[el2_ifu_mem_ctl.scala 578:57]
  reg  ifu_bus_arvalid_ff; // @[el2_ifu_mem_ctl.scala 580:53]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 592:51]
  wire  _T_2589 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 602:73]
  wire  _T_2590 = _T_2575 & _T_2589; // @[el2_ifu_mem_ctl.scala 602:71]
  wire  _T_2592 = last_data_recieved_ff & _T_1325; // @[el2_ifu_mem_ctl.scala 602:114]
  wire [2:0] _T_2598 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 607:43]
  wire  _T_2602 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 610:48]
  wire  _T_2603 = _T_2602 & miss_pending; // @[el2_ifu_mem_ctl.scala 610:68]
  wire  bus_inc_cmd_beat_cnt = _T_2603 & _T_2574; // @[el2_ifu_mem_ctl.scala 610:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 612:57]
  wire  _T_2607 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 613:31]
  wire  _T_2608 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 613:71]
  wire  _T_2609 = _T_2608 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 613:87]
  wire  _T_2610 = ~_T_2609; // @[el2_ifu_mem_ctl.scala 613:55]
  wire  bus_hold_cmd_beat_cnt = _T_2607 & _T_2610; // @[el2_ifu_mem_ctl.scala 613:53]
  wire  _T_2611 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 614:46]
  wire  bus_cmd_beat_en = _T_2611 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 614:62]
  wire [2:0] _T_2614 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 616:46]
  wire [2:0] _T_2616 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2617 = bus_inc_cmd_beat_cnt ? _T_2614 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2618 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2620 = _T_2616 | _T_2617; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2620 | _T_2618; // @[Mux.scala 27:72]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 628:62]
  wire  _T_2649 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 633:50]
  wire  _T_2650 = io_ifc_dma_access_ok & _T_2649; // @[el2_ifu_mem_ctl.scala 633:47]
  wire  _T_2651 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 633:70]
  wire  _T_2655 = _T_2650 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 634:72]
  wire  _T_2656 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 634:111]
  wire  _T_2657 = _T_2655 & _T_2656; // @[el2_ifu_mem_ctl.scala 634:97]
  wire  ifc_dma_access_q_ok = _T_2657 & _T_2651; // @[el2_ifu_mem_ctl.scala 634:127]
  wire  _T_2660 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 637:40]
  wire  _T_2661 = _T_2660 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 637:58]
  wire  _T_2664 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 638:60]
  wire  _T_2665 = _T_2660 & _T_2664; // @[el2_ifu_mem_ctl.scala 638:58]
  wire  _T_2666 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 638:104]
  wire [2:0] _T_2671 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire  _T_2692 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[33]; // @[el2_lib.scala 259:74]
  wire  _T_2693 = _T_2692 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 259:74]
  wire  _T_2694 = _T_2693 ^ io_dma_mem_wdata[36]; // @[el2_lib.scala 259:74]
  wire  _T_2695 = _T_2694 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 259:74]
  wire  _T_2696 = _T_2695 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 259:74]
  wire  _T_2697 = _T_2696 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2698 = _T_2697 ^ io_dma_mem_wdata[43]; // @[el2_lib.scala 259:74]
  wire  _T_2699 = _T_2698 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 259:74]
  wire  _T_2700 = _T_2699 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 259:74]
  wire  _T_2701 = _T_2700 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2702 = _T_2701 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 259:74]
  wire  _T_2703 = _T_2702 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2704 = _T_2703 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2705 = _T_2704 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2706 = _T_2705 ^ io_dma_mem_wdata[58]; // @[el2_lib.scala 259:74]
  wire  _T_2707 = _T_2706 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 259:74]
  wire  _T_2708 = _T_2707 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 259:74]
  wire  _T_2727 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 259:74]
  wire  _T_2728 = _T_2727 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 259:74]
  wire  _T_2729 = _T_2728 ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 259:74]
  wire  _T_2730 = _T_2729 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 259:74]
  wire  _T_2731 = _T_2730 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 259:74]
  wire  _T_2732 = _T_2731 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2733 = _T_2732 ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 259:74]
  wire  _T_2734 = _T_2733 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 259:74]
  wire  _T_2735 = _T_2734 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 259:74]
  wire  _T_2736 = _T_2735 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2737 = _T_2736 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 259:74]
  wire  _T_2738 = _T_2737 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2739 = _T_2738 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2740 = _T_2739 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2741 = _T_2740 ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 259:74]
  wire  _T_2742 = _T_2741 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 259:74]
  wire  _T_2743 = _T_2742 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 259:74]
  wire  _T_2762 = io_dma_mem_wdata[33] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 259:74]
  wire  _T_2763 = _T_2762 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 259:74]
  wire  _T_2764 = _T_2763 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 259:74]
  wire  _T_2765 = _T_2764 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 259:74]
  wire  _T_2766 = _T_2765 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 259:74]
  wire  _T_2767 = _T_2766 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2768 = _T_2767 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 259:74]
  wire  _T_2769 = _T_2768 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 259:74]
  wire  _T_2770 = _T_2769 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 259:74]
  wire  _T_2771 = _T_2770 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2772 = _T_2771 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 259:74]
  wire  _T_2773 = _T_2772 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2774 = _T_2773 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2775 = _T_2774 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2776 = _T_2775 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 259:74]
  wire  _T_2777 = _T_2776 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 259:74]
  wire  _T_2778 = _T_2777 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 259:74]
  wire  _T_2794 = io_dma_mem_wdata[36] ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 259:74]
  wire  _T_2795 = _T_2794 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 259:74]
  wire  _T_2796 = _T_2795 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 259:74]
  wire  _T_2797 = _T_2796 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 259:74]
  wire  _T_2798 = _T_2797 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 259:74]
  wire  _T_2799 = _T_2798 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2800 = _T_2799 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 259:74]
  wire  _T_2801 = _T_2800 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 259:74]
  wire  _T_2802 = _T_2801 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 259:74]
  wire  _T_2803 = _T_2802 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2804 = _T_2803 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 259:74]
  wire  _T_2805 = _T_2804 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2806 = _T_2805 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2807 = _T_2806 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2823 = io_dma_mem_wdata[43] ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 259:74]
  wire  _T_2824 = _T_2823 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 259:74]
  wire  _T_2825 = _T_2824 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 259:74]
  wire  _T_2826 = _T_2825 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 259:74]
  wire  _T_2827 = _T_2826 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 259:74]
  wire  _T_2828 = _T_2827 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2829 = _T_2828 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 259:74]
  wire  _T_2830 = _T_2829 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 259:74]
  wire  _T_2831 = _T_2830 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 259:74]
  wire  _T_2832 = _T_2831 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2833 = _T_2832 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 259:74]
  wire  _T_2834 = _T_2833 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2835 = _T_2834 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2836 = _T_2835 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2843 = io_dma_mem_wdata[58] ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 259:74]
  wire  _T_2844 = _T_2843 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 259:74]
  wire  _T_2845 = _T_2844 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 259:74]
  wire  _T_2846 = _T_2845 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 259:74]
  wire  _T_2847 = _T_2846 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 259:74]
  wire [5:0] _T_2852 = {_T_2847,_T_2836,_T_2807,_T_2778,_T_2743,_T_2708}; // @[Cat.scala 29:58]
  wire  _T_2853 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 267:13]
  wire  _T_2854 = ^_T_2852; // @[el2_lib.scala 267:23]
  wire  _T_2855 = _T_2853 ^ _T_2854; // @[el2_lib.scala 267:18]
  wire  _T_2876 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[1]; // @[el2_lib.scala 259:74]
  wire  _T_2877 = _T_2876 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 259:74]
  wire  _T_2878 = _T_2877 ^ io_dma_mem_wdata[4]; // @[el2_lib.scala 259:74]
  wire  _T_2879 = _T_2878 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 259:74]
  wire  _T_2880 = _T_2879 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 259:74]
  wire  _T_2881 = _T_2880 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_2882 = _T_2881 ^ io_dma_mem_wdata[11]; // @[el2_lib.scala 259:74]
  wire  _T_2883 = _T_2882 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 259:74]
  wire  _T_2884 = _T_2883 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 259:74]
  wire  _T_2885 = _T_2884 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_2886 = _T_2885 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 259:74]
  wire  _T_2887 = _T_2886 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_2888 = _T_2887 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_2889 = _T_2888 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_2890 = _T_2889 ^ io_dma_mem_wdata[26]; // @[el2_lib.scala 259:74]
  wire  _T_2891 = _T_2890 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 259:74]
  wire  _T_2892 = _T_2891 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 259:74]
  wire  _T_2911 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 259:74]
  wire  _T_2912 = _T_2911 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 259:74]
  wire  _T_2913 = _T_2912 ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 259:74]
  wire  _T_2914 = _T_2913 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 259:74]
  wire  _T_2915 = _T_2914 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 259:74]
  wire  _T_2916 = _T_2915 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_2917 = _T_2916 ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 259:74]
  wire  _T_2918 = _T_2917 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 259:74]
  wire  _T_2919 = _T_2918 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 259:74]
  wire  _T_2920 = _T_2919 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_2921 = _T_2920 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 259:74]
  wire  _T_2922 = _T_2921 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_2923 = _T_2922 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_2924 = _T_2923 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_2925 = _T_2924 ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 259:74]
  wire  _T_2926 = _T_2925 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 259:74]
  wire  _T_2927 = _T_2926 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 259:74]
  wire  _T_2946 = io_dma_mem_wdata[1] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 259:74]
  wire  _T_2947 = _T_2946 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 259:74]
  wire  _T_2948 = _T_2947 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 259:74]
  wire  _T_2949 = _T_2948 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 259:74]
  wire  _T_2950 = _T_2949 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 259:74]
  wire  _T_2951 = _T_2950 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_2952 = _T_2951 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 259:74]
  wire  _T_2953 = _T_2952 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 259:74]
  wire  _T_2954 = _T_2953 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 259:74]
  wire  _T_2955 = _T_2954 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_2956 = _T_2955 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 259:74]
  wire  _T_2957 = _T_2956 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_2958 = _T_2957 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_2959 = _T_2958 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_2960 = _T_2959 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 259:74]
  wire  _T_2961 = _T_2960 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 259:74]
  wire  _T_2962 = _T_2961 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 259:74]
  wire  _T_2978 = io_dma_mem_wdata[4] ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 259:74]
  wire  _T_2979 = _T_2978 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 259:74]
  wire  _T_2980 = _T_2979 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 259:74]
  wire  _T_2981 = _T_2980 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 259:74]
  wire  _T_2982 = _T_2981 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 259:74]
  wire  _T_2983 = _T_2982 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_2984 = _T_2983 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 259:74]
  wire  _T_2985 = _T_2984 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 259:74]
  wire  _T_2986 = _T_2985 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 259:74]
  wire  _T_2987 = _T_2986 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_2988 = _T_2987 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 259:74]
  wire  _T_2989 = _T_2988 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_2990 = _T_2989 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_2991 = _T_2990 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_3007 = io_dma_mem_wdata[11] ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 259:74]
  wire  _T_3008 = _T_3007 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 259:74]
  wire  _T_3009 = _T_3008 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 259:74]
  wire  _T_3010 = _T_3009 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 259:74]
  wire  _T_3011 = _T_3010 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 259:74]
  wire  _T_3012 = _T_3011 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_3013 = _T_3012 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 259:74]
  wire  _T_3014 = _T_3013 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 259:74]
  wire  _T_3015 = _T_3014 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 259:74]
  wire  _T_3016 = _T_3015 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_3017 = _T_3016 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 259:74]
  wire  _T_3018 = _T_3017 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_3019 = _T_3018 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_3020 = _T_3019 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_3027 = io_dma_mem_wdata[26] ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 259:74]
  wire  _T_3028 = _T_3027 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 259:74]
  wire  _T_3029 = _T_3028 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 259:74]
  wire  _T_3030 = _T_3029 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 259:74]
  wire  _T_3031 = _T_3030 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 259:74]
  wire [5:0] _T_3036 = {_T_3031,_T_3020,_T_2991,_T_2962,_T_2927,_T_2892}; // @[Cat.scala 29:58]
  wire  _T_3037 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 267:13]
  wire  _T_3038 = ^_T_3036; // @[el2_lib.scala 267:23]
  wire  _T_3039 = _T_3037 ^ _T_3038; // @[el2_lib.scala 267:18]
  wire [6:0] _T_3040 = {_T_3039,_T_3031,_T_3020,_T_2991,_T_2962,_T_2927,_T_2892}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2855,_T_2847,_T_2836,_T_2807,_T_2778,_T_2743,_T_2708,_T_3040}; // @[Cat.scala 29:58]
  wire  _T_3042 = ~_T_2660; // @[el2_ifu_mem_ctl.scala 644:45]
  wire  _T_3043 = iccm_correct_ecc & _T_3042; // @[el2_ifu_mem_ctl.scala 644:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3044 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3051 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 658:53]
  wire  _T_3384 = _T_3296[5:0] == 6'h27; // @[el2_lib.scala 339:41]
  wire  _T_3382 = _T_3296[5:0] == 6'h26; // @[el2_lib.scala 339:41]
  wire  _T_3380 = _T_3296[5:0] == 6'h25; // @[el2_lib.scala 339:41]
  wire  _T_3378 = _T_3296[5:0] == 6'h24; // @[el2_lib.scala 339:41]
  wire  _T_3376 = _T_3296[5:0] == 6'h23; // @[el2_lib.scala 339:41]
  wire  _T_3374 = _T_3296[5:0] == 6'h22; // @[el2_lib.scala 339:41]
  wire  _T_3372 = _T_3296[5:0] == 6'h21; // @[el2_lib.scala 339:41]
  wire  _T_3370 = _T_3296[5:0] == 6'h20; // @[el2_lib.scala 339:41]
  wire  _T_3368 = _T_3296[5:0] == 6'h1f; // @[el2_lib.scala 339:41]
  wire  _T_3366 = _T_3296[5:0] == 6'h1e; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3442 = {_T_3384,_T_3382,_T_3380,_T_3378,_T_3376,_T_3374,_T_3372,_T_3370,_T_3368,_T_3366}; // @[el2_lib.scala 342:69]
  wire  _T_3364 = _T_3296[5:0] == 6'h1d; // @[el2_lib.scala 339:41]
  wire  _T_3362 = _T_3296[5:0] == 6'h1c; // @[el2_lib.scala 339:41]
  wire  _T_3360 = _T_3296[5:0] == 6'h1b; // @[el2_lib.scala 339:41]
  wire  _T_3358 = _T_3296[5:0] == 6'h1a; // @[el2_lib.scala 339:41]
  wire  _T_3356 = _T_3296[5:0] == 6'h19; // @[el2_lib.scala 339:41]
  wire  _T_3354 = _T_3296[5:0] == 6'h18; // @[el2_lib.scala 339:41]
  wire  _T_3352 = _T_3296[5:0] == 6'h17; // @[el2_lib.scala 339:41]
  wire  _T_3350 = _T_3296[5:0] == 6'h16; // @[el2_lib.scala 339:41]
  wire  _T_3348 = _T_3296[5:0] == 6'h15; // @[el2_lib.scala 339:41]
  wire  _T_3346 = _T_3296[5:0] == 6'h14; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3433 = {_T_3364,_T_3362,_T_3360,_T_3358,_T_3356,_T_3354,_T_3352,_T_3350,_T_3348,_T_3346}; // @[el2_lib.scala 342:69]
  wire  _T_3344 = _T_3296[5:0] == 6'h13; // @[el2_lib.scala 339:41]
  wire  _T_3342 = _T_3296[5:0] == 6'h12; // @[el2_lib.scala 339:41]
  wire  _T_3340 = _T_3296[5:0] == 6'h11; // @[el2_lib.scala 339:41]
  wire  _T_3338 = _T_3296[5:0] == 6'h10; // @[el2_lib.scala 339:41]
  wire  _T_3336 = _T_3296[5:0] == 6'hf; // @[el2_lib.scala 339:41]
  wire  _T_3334 = _T_3296[5:0] == 6'he; // @[el2_lib.scala 339:41]
  wire  _T_3332 = _T_3296[5:0] == 6'hd; // @[el2_lib.scala 339:41]
  wire  _T_3330 = _T_3296[5:0] == 6'hc; // @[el2_lib.scala 339:41]
  wire  _T_3328 = _T_3296[5:0] == 6'hb; // @[el2_lib.scala 339:41]
  wire  _T_3326 = _T_3296[5:0] == 6'ha; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3423 = {_T_3344,_T_3342,_T_3340,_T_3338,_T_3336,_T_3334,_T_3332,_T_3330,_T_3328,_T_3326}; // @[el2_lib.scala 342:69]
  wire  _T_3324 = _T_3296[5:0] == 6'h9; // @[el2_lib.scala 339:41]
  wire  _T_3322 = _T_3296[5:0] == 6'h8; // @[el2_lib.scala 339:41]
  wire  _T_3320 = _T_3296[5:0] == 6'h7; // @[el2_lib.scala 339:41]
  wire  _T_3318 = _T_3296[5:0] == 6'h6; // @[el2_lib.scala 339:41]
  wire  _T_3316 = _T_3296[5:0] == 6'h5; // @[el2_lib.scala 339:41]
  wire  _T_3314 = _T_3296[5:0] == 6'h4; // @[el2_lib.scala 339:41]
  wire  _T_3312 = _T_3296[5:0] == 6'h3; // @[el2_lib.scala 339:41]
  wire  _T_3310 = _T_3296[5:0] == 6'h2; // @[el2_lib.scala 339:41]
  wire  _T_3308 = _T_3296[5:0] == 6'h1; // @[el2_lib.scala 339:41]
  wire [18:0] _T_3424 = {_T_3423,_T_3324,_T_3322,_T_3320,_T_3318,_T_3316,_T_3314,_T_3312,_T_3310,_T_3308}; // @[el2_lib.scala 342:69]
  wire [38:0] _T_3444 = {_T_3442,_T_3433,_T_3424}; // @[el2_lib.scala 342:69]
  wire [7:0] _T_3399 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3405 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3399}; // @[Cat.scala 29:58]
  wire [38:0] _T_3445 = _T_3444 ^ _T_3405; // @[el2_lib.scala 342:76]
  wire [38:0] _T_3446 = _T_3300 ? _T_3445 : _T_3405; // @[el2_lib.scala 342:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3446[37:32],_T_3446[30:16],_T_3446[14:8],_T_3446[6:4],_T_3446[2]}; // @[Cat.scala 29:58]
  wire  _T_3769 = _T_3681[5:0] == 6'h27; // @[el2_lib.scala 339:41]
  wire  _T_3767 = _T_3681[5:0] == 6'h26; // @[el2_lib.scala 339:41]
  wire  _T_3765 = _T_3681[5:0] == 6'h25; // @[el2_lib.scala 339:41]
  wire  _T_3763 = _T_3681[5:0] == 6'h24; // @[el2_lib.scala 339:41]
  wire  _T_3761 = _T_3681[5:0] == 6'h23; // @[el2_lib.scala 339:41]
  wire  _T_3759 = _T_3681[5:0] == 6'h22; // @[el2_lib.scala 339:41]
  wire  _T_3757 = _T_3681[5:0] == 6'h21; // @[el2_lib.scala 339:41]
  wire  _T_3755 = _T_3681[5:0] == 6'h20; // @[el2_lib.scala 339:41]
  wire  _T_3753 = _T_3681[5:0] == 6'h1f; // @[el2_lib.scala 339:41]
  wire  _T_3751 = _T_3681[5:0] == 6'h1e; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3827 = {_T_3769,_T_3767,_T_3765,_T_3763,_T_3761,_T_3759,_T_3757,_T_3755,_T_3753,_T_3751}; // @[el2_lib.scala 342:69]
  wire  _T_3749 = _T_3681[5:0] == 6'h1d; // @[el2_lib.scala 339:41]
  wire  _T_3747 = _T_3681[5:0] == 6'h1c; // @[el2_lib.scala 339:41]
  wire  _T_3745 = _T_3681[5:0] == 6'h1b; // @[el2_lib.scala 339:41]
  wire  _T_3743 = _T_3681[5:0] == 6'h1a; // @[el2_lib.scala 339:41]
  wire  _T_3741 = _T_3681[5:0] == 6'h19; // @[el2_lib.scala 339:41]
  wire  _T_3739 = _T_3681[5:0] == 6'h18; // @[el2_lib.scala 339:41]
  wire  _T_3737 = _T_3681[5:0] == 6'h17; // @[el2_lib.scala 339:41]
  wire  _T_3735 = _T_3681[5:0] == 6'h16; // @[el2_lib.scala 339:41]
  wire  _T_3733 = _T_3681[5:0] == 6'h15; // @[el2_lib.scala 339:41]
  wire  _T_3731 = _T_3681[5:0] == 6'h14; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3818 = {_T_3749,_T_3747,_T_3745,_T_3743,_T_3741,_T_3739,_T_3737,_T_3735,_T_3733,_T_3731}; // @[el2_lib.scala 342:69]
  wire  _T_3729 = _T_3681[5:0] == 6'h13; // @[el2_lib.scala 339:41]
  wire  _T_3727 = _T_3681[5:0] == 6'h12; // @[el2_lib.scala 339:41]
  wire  _T_3725 = _T_3681[5:0] == 6'h11; // @[el2_lib.scala 339:41]
  wire  _T_3723 = _T_3681[5:0] == 6'h10; // @[el2_lib.scala 339:41]
  wire  _T_3721 = _T_3681[5:0] == 6'hf; // @[el2_lib.scala 339:41]
  wire  _T_3719 = _T_3681[5:0] == 6'he; // @[el2_lib.scala 339:41]
  wire  _T_3717 = _T_3681[5:0] == 6'hd; // @[el2_lib.scala 339:41]
  wire  _T_3715 = _T_3681[5:0] == 6'hc; // @[el2_lib.scala 339:41]
  wire  _T_3713 = _T_3681[5:0] == 6'hb; // @[el2_lib.scala 339:41]
  wire  _T_3711 = _T_3681[5:0] == 6'ha; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3808 = {_T_3729,_T_3727,_T_3725,_T_3723,_T_3721,_T_3719,_T_3717,_T_3715,_T_3713,_T_3711}; // @[el2_lib.scala 342:69]
  wire  _T_3709 = _T_3681[5:0] == 6'h9; // @[el2_lib.scala 339:41]
  wire  _T_3707 = _T_3681[5:0] == 6'h8; // @[el2_lib.scala 339:41]
  wire  _T_3705 = _T_3681[5:0] == 6'h7; // @[el2_lib.scala 339:41]
  wire  _T_3703 = _T_3681[5:0] == 6'h6; // @[el2_lib.scala 339:41]
  wire  _T_3701 = _T_3681[5:0] == 6'h5; // @[el2_lib.scala 339:41]
  wire  _T_3699 = _T_3681[5:0] == 6'h4; // @[el2_lib.scala 339:41]
  wire  _T_3697 = _T_3681[5:0] == 6'h3; // @[el2_lib.scala 339:41]
  wire  _T_3695 = _T_3681[5:0] == 6'h2; // @[el2_lib.scala 339:41]
  wire  _T_3693 = _T_3681[5:0] == 6'h1; // @[el2_lib.scala 339:41]
  wire [18:0] _T_3809 = {_T_3808,_T_3709,_T_3707,_T_3705,_T_3703,_T_3701,_T_3699,_T_3697,_T_3695,_T_3693}; // @[el2_lib.scala 342:69]
  wire [38:0] _T_3829 = {_T_3827,_T_3818,_T_3809}; // @[el2_lib.scala 342:69]
  wire [7:0] _T_3784 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3790 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3784}; // @[Cat.scala 29:58]
  wire [38:0] _T_3830 = _T_3829 ^ _T_3790; // @[el2_lib.scala 342:76]
  wire [38:0] _T_3831 = _T_3685 ? _T_3830 : _T_3790; // @[el2_lib.scala 342:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3831[37:32],_T_3831[30:16],_T_3831[14:8],_T_3831[6:4],_T_3831[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 650:35]
  wire  _T_3304 = ~_T_3296[6]; // @[el2_lib.scala 335:55]
  wire  _T_3305 = _T_3298 & _T_3304; // @[el2_lib.scala 335:53]
  wire  _T_3689 = ~_T_3681[6]; // @[el2_lib.scala 335:55]
  wire  _T_3690 = _T_3683 & _T_3689; // @[el2_lib.scala 335:53]
  wire [1:0] iccm_double_ecc_error = {_T_3305,_T_3690}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 652:53]
  wire [63:0] _T_3055 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3056 = {iccm_dma_rdata_1_muxed,_T_3446[37:32],_T_3446[30:16],_T_3446[14:8],_T_3446[6:4],_T_3446[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 654:54]
  reg [2:0] iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 655:74]
  reg  iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 660:76]
  reg  iccm_dma_ecc_error; // @[el2_ifu_mem_ctl.scala 662:74]
  reg [63:0] iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 664:75]
  wire  _T_3061 = _T_2660 & _T_2649; // @[el2_ifu_mem_ctl.scala 667:65]
  wire  _T_3065 = _T_3042 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 668:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3066 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [14:0] _T_3068 = _T_3065 ? _T_3066 : io_ifc_fetch_addr_bf[14:0]; // @[el2_ifu_mem_ctl.scala 668:8]
  wire  _T_3458 = _T_3296 == 7'h40; // @[el2_lib.scala 345:62]
  wire  _T_3459 = _T_3446[38] ^ _T_3458; // @[el2_lib.scala 345:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3459,_T_3446[31],_T_3446[15],_T_3446[7],_T_3446[3],_T_3446[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3843 = _T_3681 == 7'h40; // @[el2_lib.scala 345:62]
  wire  _T_3844 = _T_3831[38] ^ _T_3843; // @[el2_lib.scala 345:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3844,_T_3831[31],_T_3831[15],_T_3831[7],_T_3831[3],_T_3831[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3860 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 680:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 682:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 683:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 691:62]
  wire  _T_3868 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 685:76]
  wire  _T_3869 = io_iccm_rd_ecc_single_err & _T_3868; // @[el2_ifu_mem_ctl.scala 685:74]
  wire  _T_3871 = _T_3869 & _T_319; // @[el2_ifu_mem_ctl.scala 685:104]
  wire  iccm_ecc_write_status = _T_3871 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 685:127]
  wire  _T_3872 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 686:67]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 690:51]
  wire [13:0] _T_3877 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 689:102]
  wire [38:0] _T_3881 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3886 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 694:41]
  wire  _T_3887 = io_ifc_fetch_req_bf & _T_3886; // @[el2_ifu_mem_ctl.scala 694:39]
  wire  _T_3888 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 694:72]
  wire  _T_3889 = _T_3887 & _T_3888; // @[el2_ifu_mem_ctl.scala 694:70]
  wire  _T_3891 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 695:34]
  wire  _T_3892 = _T_2219 & _T_3891; // @[el2_ifu_mem_ctl.scala 695:32]
  wire  _T_3895 = _T_2235 & _T_3891; // @[el2_ifu_mem_ctl.scala 696:37]
  wire  _T_3896 = _T_3892 | _T_3895; // @[el2_ifu_mem_ctl.scala 695:88]
  wire  _T_3897 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 697:19]
  wire  _T_3899 = _T_3897 & _T_3891; // @[el2_ifu_mem_ctl.scala 697:41]
  wire  _T_3900 = _T_3896 | _T_3899; // @[el2_ifu_mem_ctl.scala 696:88]
  wire  _T_3901 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 698:19]
  wire  _T_3903 = _T_3901 & _T_3891; // @[el2_ifu_mem_ctl.scala 698:35]
  wire  _T_3904 = _T_3900 | _T_3903; // @[el2_ifu_mem_ctl.scala 697:88]
  wire  _T_3907 = _T_2234 & _T_3891; // @[el2_ifu_mem_ctl.scala 699:38]
  wire  _T_3908 = _T_3904 | _T_3907; // @[el2_ifu_mem_ctl.scala 698:88]
  wire  _T_3910 = _T_2235 & miss_state_en; // @[el2_ifu_mem_ctl.scala 700:37]
  wire  _T_3911 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 700:71]
  wire  _T_3912 = _T_3910 & _T_3911; // @[el2_ifu_mem_ctl.scala 700:54]
  wire  _T_3913 = _T_3908 | _T_3912; // @[el2_ifu_mem_ctl.scala 699:57]
  wire  _T_3914 = ~_T_3913; // @[el2_ifu_mem_ctl.scala 695:5]
  wire  _T_3915 = _T_3889 & _T_3914; // @[el2_ifu_mem_ctl.scala 694:96]
  wire  _T_3916 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 701:26]
  wire  _T_3918 = _T_3916 & _T_3886; // @[el2_ifu_mem_ctl.scala 701:48]
  wire  _T_3920 = _T_3918 & _T_3888; // @[el2_ifu_mem_ctl.scala 701:79]
  wire [1:0] _T_3923 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9729 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 796:72]
  wire  bus_wren_1 = _T_9729 & miss_pending; // @[el2_ifu_mem_ctl.scala 796:96]
  wire  _T_9728 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 796:72]
  wire  bus_wren_0 = _T_9728 & miss_pending; // @[el2_ifu_mem_ctl.scala 796:96]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_3929 = ~_T_108; // @[el2_ifu_mem_ctl.scala 704:106]
  wire  _T_3930 = _T_2219 & _T_3929; // @[el2_ifu_mem_ctl.scala 704:104]
  wire  _T_3931 = _T_2235 | _T_3930; // @[el2_ifu_mem_ctl.scala 704:77]
  wire  _T_3935 = ~_T_51; // @[el2_ifu_mem_ctl.scala 704:172]
  wire  _T_3936 = _T_3931 & _T_3935; // @[el2_ifu_mem_ctl.scala 704:170]
  wire  _T_3937 = ~_T_3936; // @[el2_ifu_mem_ctl.scala 704:44]
  wire  _T_3941 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 707:62]
  wire  _T_3942 = ~_T_3941; // @[el2_ifu_mem_ctl.scala 707:48]
  wire  _T_3943 = _T_276 & _T_3942; // @[el2_ifu_mem_ctl.scala 707:46]
  wire  _T_3944 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 707:79]
  wire  ic_valid = _T_3943 & _T_3944; // @[el2_ifu_mem_ctl.scala 707:77]
  wire  _T_3946 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 708:80]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 711:12]
  wire  _T_3949 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 714:72]
  wire  _T_9726 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 795:43]
  wire  way_status_wr_en = _T_9726 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 795:56]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 716:12]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 791:39]
  reg  way_status_new_ff; // @[el2_ifu_mem_ctl.scala 722:12]
  wire  _T_3969 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[el2_ifu_mem_ctl.scala 728:126]
  wire  _T_3970 = _T_3969 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:134]
  wire  _T_3973 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[el2_ifu_mem_ctl.scala 728:126]
  wire  _T_3974 = _T_3973 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:134]
  wire  _T_3977 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[el2_ifu_mem_ctl.scala 728:126]
  wire  _T_3978 = _T_3977 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:134]
  wire  _T_3981 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[el2_ifu_mem_ctl.scala 728:126]
  wire  _T_3982 = _T_3981 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:134]
  wire  _T_3985 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[el2_ifu_mem_ctl.scala 728:126]
  wire  _T_3986 = _T_3985 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:134]
  wire  _T_3989 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[el2_ifu_mem_ctl.scala 728:126]
  wire  _T_3990 = _T_3989 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:134]
  wire  _T_3993 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[el2_ifu_mem_ctl.scala 728:126]
  wire  _T_3994 = _T_3993 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:134]
  wire  _T_3997 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[el2_ifu_mem_ctl.scala 728:126]
  wire  _T_3998 = _T_3997 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:134]
  wire  _T_9732 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 798:82]
  wire  _T_9733 = _T_9732 & miss_pending; // @[el2_ifu_mem_ctl.scala 798:106]
  wire  bus_wren_last_1 = _T_9733 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 798:121]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 799:82]
  wire  _T_9735 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 800:71]
  wire  _T_9730 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 798:82]
  wire  _T_9731 = _T_9730 & miss_pending; // @[el2_ifu_mem_ctl.scala 798:106]
  wire  bus_wren_last_0 = _T_9731 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 798:121]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 799:82]
  wire  _T_9734 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 800:71]
  wire [1:0] ifu_tag_wren = {_T_9735,_T_9734}; // @[Cat.scala 29:58]
  wire [1:0] _T_9770 = _T_3949 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9770 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 834:90]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 743:12]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 747:12]
  wire  _T_5012 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 751:76]
  wire  _T_5014 = _T_5012 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:85]
  wire  _T_5016 = perr_ic_index_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 752:68]
  wire  _T_5018 = _T_5016 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 752:77]
  wire  _T_5019 = _T_5014 | _T_5018; // @[el2_ifu_mem_ctl.scala 751:107]
  wire  _T_5020 = _T_5019 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:100]
  wire  _T_5024 = _T_5012 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:85]
  wire  _T_5028 = _T_5016 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 752:77]
  wire  _T_5029 = _T_5024 | _T_5028; // @[el2_ifu_mem_ctl.scala 751:107]
  wire  _T_5030 = _T_5029 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:100]
  wire [1:0] tag_valid_clken_0 = {_T_5030,_T_5020}; // @[Cat.scala 29:58]
  wire  _T_5032 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 751:76]
  wire  _T_5034 = _T_5032 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:85]
  wire  _T_5036 = perr_ic_index_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 752:68]
  wire  _T_5038 = _T_5036 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 752:77]
  wire  _T_5039 = _T_5034 | _T_5038; // @[el2_ifu_mem_ctl.scala 751:107]
  wire  _T_5040 = _T_5039 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:100]
  wire  _T_5044 = _T_5032 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:85]
  wire  _T_5048 = _T_5036 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 752:77]
  wire  _T_5049 = _T_5044 | _T_5048; // @[el2_ifu_mem_ctl.scala 751:107]
  wire  _T_5050 = _T_5049 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:100]
  wire [1:0] tag_valid_clken_1 = {_T_5050,_T_5040}; // @[Cat.scala 29:58]
  wire  _T_5052 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 751:76]
  wire  _T_5054 = _T_5052 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:85]
  wire  _T_5056 = perr_ic_index_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 752:68]
  wire  _T_5058 = _T_5056 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 752:77]
  wire  _T_5059 = _T_5054 | _T_5058; // @[el2_ifu_mem_ctl.scala 751:107]
  wire  _T_5060 = _T_5059 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:100]
  wire  _T_5064 = _T_5052 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:85]
  wire  _T_5068 = _T_5056 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 752:77]
  wire  _T_5069 = _T_5064 | _T_5068; // @[el2_ifu_mem_ctl.scala 751:107]
  wire  _T_5070 = _T_5069 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:100]
  wire [1:0] tag_valid_clken_2 = {_T_5070,_T_5060}; // @[Cat.scala 29:58]
  wire  _T_5072 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 751:76]
  wire  _T_5074 = _T_5072 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:85]
  wire  _T_5076 = perr_ic_index_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 752:68]
  wire  _T_5078 = _T_5076 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 752:77]
  wire  _T_5079 = _T_5074 | _T_5078; // @[el2_ifu_mem_ctl.scala 751:107]
  wire  _T_5080 = _T_5079 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:100]
  wire  _T_5084 = _T_5072 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:85]
  wire  _T_5088 = _T_5076 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 752:77]
  wire  _T_5089 = _T_5084 | _T_5088; // @[el2_ifu_mem_ctl.scala 751:107]
  wire  _T_5090 = _T_5089 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:100]
  wire [1:0] tag_valid_clken_3 = {_T_5090,_T_5080}; // @[Cat.scala 29:58]
  wire  _T_5101 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 760:95]
  wire  _T_5102 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 760:122]
  wire  _T_5103 = _T_5101 & _T_5102; // @[el2_ifu_mem_ctl.scala 760:120]
  wire  _T_5106 = _T_4620 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5107 = perr_ic_index_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5109 = _T_5107 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5110 = _T_5106 | _T_5109; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5111 = _T_5110 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5121 = _T_4621 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5122 = perr_ic_index_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5124 = _T_5122 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5125 = _T_5121 | _T_5124; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5126 = _T_5125 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5136 = _T_4622 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5137 = perr_ic_index_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5139 = _T_5137 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5140 = _T_5136 | _T_5139; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5141 = _T_5140 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5151 = _T_4623 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5152 = perr_ic_index_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5154 = _T_5152 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5155 = _T_5151 | _T_5154; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5156 = _T_5155 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5166 = _T_4624 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5167 = perr_ic_index_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5169 = _T_5167 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5170 = _T_5166 | _T_5169; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5171 = _T_5170 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5181 = _T_4625 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5182 = perr_ic_index_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5184 = _T_5182 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5185 = _T_5181 | _T_5184; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5186 = _T_5185 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5196 = _T_4626 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5197 = perr_ic_index_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5199 = _T_5197 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5200 = _T_5196 | _T_5199; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5201 = _T_5200 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5211 = _T_4627 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5212 = perr_ic_index_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5214 = _T_5212 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5215 = _T_5211 | _T_5214; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5216 = _T_5215 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5226 = _T_4628 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5227 = perr_ic_index_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5229 = _T_5227 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5230 = _T_5226 | _T_5229; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5231 = _T_5230 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5241 = _T_4629 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5242 = perr_ic_index_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5244 = _T_5242 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5245 = _T_5241 | _T_5244; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5246 = _T_5245 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5256 = _T_4630 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5257 = perr_ic_index_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5259 = _T_5257 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5260 = _T_5256 | _T_5259; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5261 = _T_5260 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5271 = _T_4631 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5272 = perr_ic_index_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5274 = _T_5272 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5275 = _T_5271 | _T_5274; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5276 = _T_5275 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5286 = _T_4632 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5287 = perr_ic_index_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5289 = _T_5287 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5290 = _T_5286 | _T_5289; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5291 = _T_5290 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5301 = _T_4633 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5302 = perr_ic_index_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5304 = _T_5302 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5305 = _T_5301 | _T_5304; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5306 = _T_5305 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5316 = _T_4634 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5317 = perr_ic_index_ff == 7'he; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5319 = _T_5317 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5320 = _T_5316 | _T_5319; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5321 = _T_5320 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5331 = _T_4635 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5332 = perr_ic_index_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5334 = _T_5332 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5335 = _T_5331 | _T_5334; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5336 = _T_5335 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5346 = _T_4636 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5347 = perr_ic_index_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5349 = _T_5347 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5350 = _T_5346 | _T_5349; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5351 = _T_5350 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5361 = _T_4637 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5362 = perr_ic_index_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5364 = _T_5362 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5365 = _T_5361 | _T_5364; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5366 = _T_5365 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5376 = _T_4638 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5377 = perr_ic_index_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5379 = _T_5377 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5380 = _T_5376 | _T_5379; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5381 = _T_5380 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5391 = _T_4639 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5392 = perr_ic_index_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5394 = _T_5392 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5395 = _T_5391 | _T_5394; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5396 = _T_5395 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5406 = _T_4640 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5407 = perr_ic_index_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5409 = _T_5407 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5410 = _T_5406 | _T_5409; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5411 = _T_5410 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5421 = _T_4641 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5422 = perr_ic_index_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5424 = _T_5422 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5425 = _T_5421 | _T_5424; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5426 = _T_5425 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5436 = _T_4642 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5437 = perr_ic_index_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5439 = _T_5437 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5440 = _T_5436 | _T_5439; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5441 = _T_5440 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5451 = _T_4643 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5452 = perr_ic_index_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5454 = _T_5452 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5455 = _T_5451 | _T_5454; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5456 = _T_5455 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5466 = _T_4644 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5467 = perr_ic_index_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5469 = _T_5467 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5470 = _T_5466 | _T_5469; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5471 = _T_5470 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5481 = _T_4645 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5482 = perr_ic_index_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5484 = _T_5482 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5485 = _T_5481 | _T_5484; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5486 = _T_5485 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5496 = _T_4646 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5497 = perr_ic_index_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5499 = _T_5497 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5500 = _T_5496 | _T_5499; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5501 = _T_5500 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5511 = _T_4647 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5512 = perr_ic_index_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5514 = _T_5512 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5515 = _T_5511 | _T_5514; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5516 = _T_5515 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5526 = _T_4648 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5527 = perr_ic_index_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5529 = _T_5527 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5530 = _T_5526 | _T_5529; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5531 = _T_5530 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5541 = _T_4649 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5542 = perr_ic_index_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5544 = _T_5542 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5545 = _T_5541 | _T_5544; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5546 = _T_5545 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5556 = _T_4650 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5557 = perr_ic_index_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5559 = _T_5557 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5560 = _T_5556 | _T_5559; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5561 = _T_5560 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5571 = _T_4651 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5572 = perr_ic_index_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_5574 = _T_5572 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5575 = _T_5571 | _T_5574; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5576 = _T_5575 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5586 = _T_4620 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5589 = _T_5107 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5590 = _T_5586 | _T_5589; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5591 = _T_5590 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5601 = _T_4621 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5604 = _T_5122 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5605 = _T_5601 | _T_5604; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5606 = _T_5605 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5616 = _T_4622 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5619 = _T_5137 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5620 = _T_5616 | _T_5619; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5621 = _T_5620 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5631 = _T_4623 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5634 = _T_5152 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5635 = _T_5631 | _T_5634; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5636 = _T_5635 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5646 = _T_4624 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5649 = _T_5167 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5650 = _T_5646 | _T_5649; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5651 = _T_5650 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5661 = _T_4625 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5664 = _T_5182 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5665 = _T_5661 | _T_5664; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5666 = _T_5665 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5676 = _T_4626 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5679 = _T_5197 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5680 = _T_5676 | _T_5679; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5681 = _T_5680 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5691 = _T_4627 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5694 = _T_5212 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5695 = _T_5691 | _T_5694; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5696 = _T_5695 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5706 = _T_4628 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5709 = _T_5227 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5710 = _T_5706 | _T_5709; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5711 = _T_5710 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5721 = _T_4629 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5724 = _T_5242 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5725 = _T_5721 | _T_5724; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5726 = _T_5725 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5736 = _T_4630 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5739 = _T_5257 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5740 = _T_5736 | _T_5739; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5741 = _T_5740 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5751 = _T_4631 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5754 = _T_5272 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5755 = _T_5751 | _T_5754; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5756 = _T_5755 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5766 = _T_4632 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5769 = _T_5287 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5770 = _T_5766 | _T_5769; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5771 = _T_5770 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5781 = _T_4633 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5784 = _T_5302 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5785 = _T_5781 | _T_5784; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5786 = _T_5785 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5796 = _T_4634 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5799 = _T_5317 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5800 = _T_5796 | _T_5799; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5801 = _T_5800 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5811 = _T_4635 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5814 = _T_5332 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5815 = _T_5811 | _T_5814; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5816 = _T_5815 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5826 = _T_4636 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5829 = _T_5347 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5830 = _T_5826 | _T_5829; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5831 = _T_5830 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5841 = _T_4637 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5844 = _T_5362 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5845 = _T_5841 | _T_5844; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5846 = _T_5845 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5856 = _T_4638 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5859 = _T_5377 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5860 = _T_5856 | _T_5859; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5861 = _T_5860 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5871 = _T_4639 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5874 = _T_5392 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5875 = _T_5871 | _T_5874; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5876 = _T_5875 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5886 = _T_4640 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5889 = _T_5407 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5890 = _T_5886 | _T_5889; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5891 = _T_5890 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5901 = _T_4641 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5904 = _T_5422 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5905 = _T_5901 | _T_5904; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5906 = _T_5905 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5916 = _T_4642 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5919 = _T_5437 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5920 = _T_5916 | _T_5919; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5921 = _T_5920 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5931 = _T_4643 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5934 = _T_5452 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5935 = _T_5931 | _T_5934; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5936 = _T_5935 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5946 = _T_4644 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5949 = _T_5467 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5950 = _T_5946 | _T_5949; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5951 = _T_5950 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5961 = _T_4645 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5964 = _T_5482 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5965 = _T_5961 | _T_5964; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5966 = _T_5965 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5976 = _T_4646 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5979 = _T_5497 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5980 = _T_5976 | _T_5979; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5981 = _T_5980 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_5991 = _T_4647 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_5994 = _T_5512 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_5995 = _T_5991 | _T_5994; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_5996 = _T_5995 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6006 = _T_4648 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6009 = _T_5527 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6010 = _T_6006 | _T_6009; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6011 = _T_6010 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6021 = _T_4649 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6024 = _T_5542 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6025 = _T_6021 | _T_6024; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6026 = _T_6025 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6036 = _T_4650 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6039 = _T_5557 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6040 = _T_6036 | _T_6039; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6041 = _T_6040 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6051 = _T_4651 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6054 = _T_5572 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6055 = _T_6051 | _T_6054; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6056 = _T_6055 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6066 = _T_4652 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6067 = perr_ic_index_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6069 = _T_6067 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6070 = _T_6066 | _T_6069; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6071 = _T_6070 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6081 = _T_4653 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6082 = perr_ic_index_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6084 = _T_6082 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6085 = _T_6081 | _T_6084; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6086 = _T_6085 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6096 = _T_4654 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6097 = perr_ic_index_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6099 = _T_6097 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6100 = _T_6096 | _T_6099; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6101 = _T_6100 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6111 = _T_4655 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6112 = perr_ic_index_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6114 = _T_6112 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6115 = _T_6111 | _T_6114; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6116 = _T_6115 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6126 = _T_4656 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6127 = perr_ic_index_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6129 = _T_6127 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6130 = _T_6126 | _T_6129; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6131 = _T_6130 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6141 = _T_4657 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6142 = perr_ic_index_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6144 = _T_6142 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6145 = _T_6141 | _T_6144; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6146 = _T_6145 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6156 = _T_4658 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6157 = perr_ic_index_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6159 = _T_6157 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6160 = _T_6156 | _T_6159; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6161 = _T_6160 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6171 = _T_4659 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6172 = perr_ic_index_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6174 = _T_6172 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6175 = _T_6171 | _T_6174; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6176 = _T_6175 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6186 = _T_4660 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6187 = perr_ic_index_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6189 = _T_6187 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6190 = _T_6186 | _T_6189; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6191 = _T_6190 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6201 = _T_4661 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6202 = perr_ic_index_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6204 = _T_6202 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6205 = _T_6201 | _T_6204; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6206 = _T_6205 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6216 = _T_4662 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6217 = perr_ic_index_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6219 = _T_6217 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6220 = _T_6216 | _T_6219; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6221 = _T_6220 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6231 = _T_4663 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6232 = perr_ic_index_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6234 = _T_6232 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6235 = _T_6231 | _T_6234; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6236 = _T_6235 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6246 = _T_4664 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6247 = perr_ic_index_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6249 = _T_6247 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6250 = _T_6246 | _T_6249; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6251 = _T_6250 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6261 = _T_4665 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6262 = perr_ic_index_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6264 = _T_6262 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6265 = _T_6261 | _T_6264; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6266 = _T_6265 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6276 = _T_4666 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6277 = perr_ic_index_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6279 = _T_6277 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6280 = _T_6276 | _T_6279; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6281 = _T_6280 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6291 = _T_4667 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6292 = perr_ic_index_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6294 = _T_6292 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6295 = _T_6291 | _T_6294; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6296 = _T_6295 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6306 = _T_4668 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6307 = perr_ic_index_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6309 = _T_6307 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6310 = _T_6306 | _T_6309; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6311 = _T_6310 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6321 = _T_4669 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6322 = perr_ic_index_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6324 = _T_6322 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6325 = _T_6321 | _T_6324; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6326 = _T_6325 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6336 = _T_4670 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6337 = perr_ic_index_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6339 = _T_6337 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6340 = _T_6336 | _T_6339; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6341 = _T_6340 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6351 = _T_4671 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6352 = perr_ic_index_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6354 = _T_6352 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6355 = _T_6351 | _T_6354; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6356 = _T_6355 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6366 = _T_4672 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6367 = perr_ic_index_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6369 = _T_6367 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6370 = _T_6366 | _T_6369; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6371 = _T_6370 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6381 = _T_4673 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6382 = perr_ic_index_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6384 = _T_6382 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6385 = _T_6381 | _T_6384; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6386 = _T_6385 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6396 = _T_4674 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6397 = perr_ic_index_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6399 = _T_6397 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6400 = _T_6396 | _T_6399; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6401 = _T_6400 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6411 = _T_4675 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6412 = perr_ic_index_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6414 = _T_6412 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6415 = _T_6411 | _T_6414; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6416 = _T_6415 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6426 = _T_4676 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6427 = perr_ic_index_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6429 = _T_6427 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6430 = _T_6426 | _T_6429; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6431 = _T_6430 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6441 = _T_4677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6442 = perr_ic_index_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6444 = _T_6442 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6445 = _T_6441 | _T_6444; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6446 = _T_6445 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6456 = _T_4678 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6457 = perr_ic_index_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6459 = _T_6457 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6460 = _T_6456 | _T_6459; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6461 = _T_6460 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6471 = _T_4679 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6472 = perr_ic_index_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6474 = _T_6472 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6475 = _T_6471 | _T_6474; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6476 = _T_6475 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6486 = _T_4680 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6487 = perr_ic_index_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6489 = _T_6487 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6490 = _T_6486 | _T_6489; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6491 = _T_6490 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6501 = _T_4681 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6502 = perr_ic_index_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6504 = _T_6502 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6505 = _T_6501 | _T_6504; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6506 = _T_6505 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6516 = _T_4682 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6517 = perr_ic_index_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6519 = _T_6517 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6520 = _T_6516 | _T_6519; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6521 = _T_6520 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6531 = _T_4683 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6532 = perr_ic_index_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_6534 = _T_6532 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6535 = _T_6531 | _T_6534; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6536 = _T_6535 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6546 = _T_4652 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6549 = _T_6067 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6550 = _T_6546 | _T_6549; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6551 = _T_6550 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6561 = _T_4653 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6564 = _T_6082 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6565 = _T_6561 | _T_6564; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6566 = _T_6565 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6576 = _T_4654 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6579 = _T_6097 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6580 = _T_6576 | _T_6579; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6581 = _T_6580 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6591 = _T_4655 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6594 = _T_6112 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6595 = _T_6591 | _T_6594; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6596 = _T_6595 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6606 = _T_4656 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6609 = _T_6127 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6610 = _T_6606 | _T_6609; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6611 = _T_6610 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6621 = _T_4657 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6624 = _T_6142 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6625 = _T_6621 | _T_6624; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6626 = _T_6625 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6636 = _T_4658 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6639 = _T_6157 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6640 = _T_6636 | _T_6639; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6641 = _T_6640 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6651 = _T_4659 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6654 = _T_6172 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6655 = _T_6651 | _T_6654; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6656 = _T_6655 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6666 = _T_4660 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6669 = _T_6187 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6670 = _T_6666 | _T_6669; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6671 = _T_6670 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6681 = _T_4661 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6684 = _T_6202 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6685 = _T_6681 | _T_6684; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6686 = _T_6685 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6696 = _T_4662 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6699 = _T_6217 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6700 = _T_6696 | _T_6699; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6701 = _T_6700 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6711 = _T_4663 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6714 = _T_6232 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6715 = _T_6711 | _T_6714; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6716 = _T_6715 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6726 = _T_4664 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6729 = _T_6247 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6730 = _T_6726 | _T_6729; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6731 = _T_6730 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6741 = _T_4665 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6744 = _T_6262 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6745 = _T_6741 | _T_6744; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6746 = _T_6745 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6756 = _T_4666 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6759 = _T_6277 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6760 = _T_6756 | _T_6759; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6761 = _T_6760 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6771 = _T_4667 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6774 = _T_6292 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6775 = _T_6771 | _T_6774; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6776 = _T_6775 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6786 = _T_4668 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6789 = _T_6307 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6790 = _T_6786 | _T_6789; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6791 = _T_6790 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6801 = _T_4669 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6804 = _T_6322 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6805 = _T_6801 | _T_6804; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6806 = _T_6805 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6816 = _T_4670 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6819 = _T_6337 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6820 = _T_6816 | _T_6819; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6821 = _T_6820 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6831 = _T_4671 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6834 = _T_6352 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6835 = _T_6831 | _T_6834; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6836 = _T_6835 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6846 = _T_4672 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6849 = _T_6367 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6850 = _T_6846 | _T_6849; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6851 = _T_6850 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6861 = _T_4673 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6864 = _T_6382 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6865 = _T_6861 | _T_6864; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6866 = _T_6865 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6876 = _T_4674 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6879 = _T_6397 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6880 = _T_6876 | _T_6879; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6881 = _T_6880 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6891 = _T_4675 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6894 = _T_6412 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6895 = _T_6891 | _T_6894; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6896 = _T_6895 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6906 = _T_4676 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6909 = _T_6427 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6910 = _T_6906 | _T_6909; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6911 = _T_6910 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6921 = _T_4677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6924 = _T_6442 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6925 = _T_6921 | _T_6924; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6926 = _T_6925 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6936 = _T_4678 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6939 = _T_6457 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6940 = _T_6936 | _T_6939; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6941 = _T_6940 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6951 = _T_4679 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6954 = _T_6472 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6955 = _T_6951 | _T_6954; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6956 = _T_6955 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6966 = _T_4680 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6969 = _T_6487 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6970 = _T_6966 | _T_6969; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6971 = _T_6970 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6981 = _T_4681 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6984 = _T_6502 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_6985 = _T_6981 | _T_6984; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_6986 = _T_6985 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_6996 = _T_4682 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_6999 = _T_6517 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7000 = _T_6996 | _T_6999; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7001 = _T_7000 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7011 = _T_4683 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7014 = _T_6532 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7015 = _T_7011 | _T_7014; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7016 = _T_7015 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7026 = _T_4684 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7027 = perr_ic_index_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7029 = _T_7027 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7030 = _T_7026 | _T_7029; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7031 = _T_7030 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7041 = _T_4685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7042 = perr_ic_index_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7044 = _T_7042 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7045 = _T_7041 | _T_7044; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7046 = _T_7045 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7056 = _T_4686 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7057 = perr_ic_index_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7059 = _T_7057 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7060 = _T_7056 | _T_7059; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7061 = _T_7060 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7071 = _T_4687 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7072 = perr_ic_index_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7074 = _T_7072 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7075 = _T_7071 | _T_7074; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7076 = _T_7075 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7086 = _T_4688 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7087 = perr_ic_index_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7089 = _T_7087 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7090 = _T_7086 | _T_7089; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7091 = _T_7090 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7101 = _T_4689 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7102 = perr_ic_index_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7104 = _T_7102 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7105 = _T_7101 | _T_7104; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7106 = _T_7105 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7116 = _T_4690 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7117 = perr_ic_index_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7119 = _T_7117 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7120 = _T_7116 | _T_7119; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7121 = _T_7120 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7131 = _T_4691 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7132 = perr_ic_index_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7134 = _T_7132 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7135 = _T_7131 | _T_7134; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7136 = _T_7135 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7146 = _T_4692 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7147 = perr_ic_index_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7149 = _T_7147 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7150 = _T_7146 | _T_7149; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7151 = _T_7150 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7161 = _T_4693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7162 = perr_ic_index_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7164 = _T_7162 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7165 = _T_7161 | _T_7164; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7166 = _T_7165 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7176 = _T_4694 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7177 = perr_ic_index_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7179 = _T_7177 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7180 = _T_7176 | _T_7179; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7181 = _T_7180 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7191 = _T_4695 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7192 = perr_ic_index_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7194 = _T_7192 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7195 = _T_7191 | _T_7194; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7196 = _T_7195 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7206 = _T_4696 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7207 = perr_ic_index_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7209 = _T_7207 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7210 = _T_7206 | _T_7209; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7211 = _T_7210 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7221 = _T_4697 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7222 = perr_ic_index_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7224 = _T_7222 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7225 = _T_7221 | _T_7224; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7226 = _T_7225 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7236 = _T_4698 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7237 = perr_ic_index_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7239 = _T_7237 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7240 = _T_7236 | _T_7239; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7241 = _T_7240 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7251 = _T_4699 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7252 = perr_ic_index_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7254 = _T_7252 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7255 = _T_7251 | _T_7254; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7256 = _T_7255 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7266 = _T_4700 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7267 = perr_ic_index_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7269 = _T_7267 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7270 = _T_7266 | _T_7269; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7271 = _T_7270 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7281 = _T_4701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7282 = perr_ic_index_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7284 = _T_7282 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7285 = _T_7281 | _T_7284; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7286 = _T_7285 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7296 = _T_4702 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7297 = perr_ic_index_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7299 = _T_7297 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7300 = _T_7296 | _T_7299; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7301 = _T_7300 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7311 = _T_4703 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7312 = perr_ic_index_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7314 = _T_7312 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7315 = _T_7311 | _T_7314; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7316 = _T_7315 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7326 = _T_4704 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7327 = perr_ic_index_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7329 = _T_7327 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7330 = _T_7326 | _T_7329; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7331 = _T_7330 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7341 = _T_4705 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7342 = perr_ic_index_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7344 = _T_7342 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7345 = _T_7341 | _T_7344; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7346 = _T_7345 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7356 = _T_4706 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7357 = perr_ic_index_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7359 = _T_7357 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7360 = _T_7356 | _T_7359; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7361 = _T_7360 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7371 = _T_4707 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7372 = perr_ic_index_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7374 = _T_7372 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7375 = _T_7371 | _T_7374; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7376 = _T_7375 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7386 = _T_4708 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7387 = perr_ic_index_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7389 = _T_7387 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7390 = _T_7386 | _T_7389; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7391 = _T_7390 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7401 = _T_4709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7402 = perr_ic_index_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7404 = _T_7402 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7405 = _T_7401 | _T_7404; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7406 = _T_7405 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7416 = _T_4710 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7417 = perr_ic_index_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7419 = _T_7417 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7420 = _T_7416 | _T_7419; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7421 = _T_7420 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7431 = _T_4711 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7432 = perr_ic_index_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7434 = _T_7432 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7435 = _T_7431 | _T_7434; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7436 = _T_7435 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7446 = _T_4712 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7447 = perr_ic_index_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7449 = _T_7447 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7450 = _T_7446 | _T_7449; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7451 = _T_7450 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7461 = _T_4713 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7462 = perr_ic_index_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7464 = _T_7462 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7465 = _T_7461 | _T_7464; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7466 = _T_7465 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7476 = _T_4714 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7477 = perr_ic_index_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7479 = _T_7477 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7480 = _T_7476 | _T_7479; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7481 = _T_7480 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7491 = _T_4715 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7492 = perr_ic_index_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7494 = _T_7492 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7495 = _T_7491 | _T_7494; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7496 = _T_7495 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7506 = _T_4684 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7509 = _T_7027 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7510 = _T_7506 | _T_7509; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7511 = _T_7510 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7521 = _T_4685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7524 = _T_7042 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7525 = _T_7521 | _T_7524; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7526 = _T_7525 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7536 = _T_4686 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7539 = _T_7057 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7540 = _T_7536 | _T_7539; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7541 = _T_7540 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7551 = _T_4687 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7554 = _T_7072 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7555 = _T_7551 | _T_7554; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7556 = _T_7555 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7566 = _T_4688 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7569 = _T_7087 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7570 = _T_7566 | _T_7569; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7571 = _T_7570 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7581 = _T_4689 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7584 = _T_7102 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7585 = _T_7581 | _T_7584; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7586 = _T_7585 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7596 = _T_4690 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7599 = _T_7117 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7600 = _T_7596 | _T_7599; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7601 = _T_7600 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7611 = _T_4691 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7614 = _T_7132 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7615 = _T_7611 | _T_7614; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7616 = _T_7615 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7626 = _T_4692 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7629 = _T_7147 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7630 = _T_7626 | _T_7629; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7631 = _T_7630 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7641 = _T_4693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7644 = _T_7162 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7645 = _T_7641 | _T_7644; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7646 = _T_7645 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7656 = _T_4694 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7659 = _T_7177 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7660 = _T_7656 | _T_7659; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7661 = _T_7660 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7671 = _T_4695 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7674 = _T_7192 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7675 = _T_7671 | _T_7674; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7676 = _T_7675 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7686 = _T_4696 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7689 = _T_7207 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7690 = _T_7686 | _T_7689; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7691 = _T_7690 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7701 = _T_4697 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7704 = _T_7222 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7705 = _T_7701 | _T_7704; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7706 = _T_7705 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7716 = _T_4698 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7719 = _T_7237 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7720 = _T_7716 | _T_7719; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7721 = _T_7720 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7731 = _T_4699 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7734 = _T_7252 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7735 = _T_7731 | _T_7734; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7736 = _T_7735 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7746 = _T_4700 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7749 = _T_7267 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7750 = _T_7746 | _T_7749; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7751 = _T_7750 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7761 = _T_4701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7764 = _T_7282 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7765 = _T_7761 | _T_7764; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7766 = _T_7765 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7776 = _T_4702 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7779 = _T_7297 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7780 = _T_7776 | _T_7779; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7781 = _T_7780 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7791 = _T_4703 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7794 = _T_7312 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7795 = _T_7791 | _T_7794; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7796 = _T_7795 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7806 = _T_4704 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7809 = _T_7327 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7810 = _T_7806 | _T_7809; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7811 = _T_7810 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7821 = _T_4705 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7824 = _T_7342 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7825 = _T_7821 | _T_7824; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7826 = _T_7825 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7836 = _T_4706 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7839 = _T_7357 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7840 = _T_7836 | _T_7839; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7841 = _T_7840 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7851 = _T_4707 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7854 = _T_7372 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7855 = _T_7851 | _T_7854; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7856 = _T_7855 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7866 = _T_4708 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7869 = _T_7387 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7870 = _T_7866 | _T_7869; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7871 = _T_7870 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7881 = _T_4709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7884 = _T_7402 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7885 = _T_7881 | _T_7884; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7886 = _T_7885 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7896 = _T_4710 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7899 = _T_7417 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7900 = _T_7896 | _T_7899; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7901 = _T_7900 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7911 = _T_4711 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7914 = _T_7432 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7915 = _T_7911 | _T_7914; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7916 = _T_7915 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7926 = _T_4712 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7929 = _T_7447 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7930 = _T_7926 | _T_7929; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7931 = _T_7930 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7941 = _T_4713 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7944 = _T_7462 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7945 = _T_7941 | _T_7944; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7946 = _T_7945 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7956 = _T_4714 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7959 = _T_7477 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7960 = _T_7956 | _T_7959; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7961 = _T_7960 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7971 = _T_4715 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7974 = _T_7492 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7975 = _T_7971 | _T_7974; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7976 = _T_7975 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_7986 = _T_4716 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_7987 = perr_ic_index_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_7989 = _T_7987 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_7990 = _T_7986 | _T_7989; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_7991 = _T_7990 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8001 = _T_4717 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8002 = perr_ic_index_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8004 = _T_8002 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8005 = _T_8001 | _T_8004; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8006 = _T_8005 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8016 = _T_4718 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8017 = perr_ic_index_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8019 = _T_8017 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8020 = _T_8016 | _T_8019; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8021 = _T_8020 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8031 = _T_4719 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8032 = perr_ic_index_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8034 = _T_8032 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8035 = _T_8031 | _T_8034; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8036 = _T_8035 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8046 = _T_4720 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8047 = perr_ic_index_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8049 = _T_8047 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8050 = _T_8046 | _T_8049; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8051 = _T_8050 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8061 = _T_4721 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8062 = perr_ic_index_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8064 = _T_8062 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8065 = _T_8061 | _T_8064; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8066 = _T_8065 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8076 = _T_4722 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8077 = perr_ic_index_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8079 = _T_8077 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8080 = _T_8076 | _T_8079; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8081 = _T_8080 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8091 = _T_4723 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8092 = perr_ic_index_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8094 = _T_8092 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8095 = _T_8091 | _T_8094; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8096 = _T_8095 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8106 = _T_4724 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8107 = perr_ic_index_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8109 = _T_8107 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8110 = _T_8106 | _T_8109; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8111 = _T_8110 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8121 = _T_4725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8122 = perr_ic_index_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8124 = _T_8122 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8125 = _T_8121 | _T_8124; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8126 = _T_8125 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8136 = _T_4726 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8137 = perr_ic_index_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8139 = _T_8137 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8140 = _T_8136 | _T_8139; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8141 = _T_8140 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8151 = _T_4727 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8152 = perr_ic_index_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8154 = _T_8152 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8155 = _T_8151 | _T_8154; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8156 = _T_8155 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8166 = _T_4728 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8167 = perr_ic_index_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8169 = _T_8167 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8170 = _T_8166 | _T_8169; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8171 = _T_8170 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8181 = _T_4729 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8182 = perr_ic_index_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8184 = _T_8182 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8185 = _T_8181 | _T_8184; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8186 = _T_8185 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8196 = _T_4730 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8197 = perr_ic_index_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8199 = _T_8197 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8200 = _T_8196 | _T_8199; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8201 = _T_8200 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8211 = _T_4731 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8212 = perr_ic_index_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8214 = _T_8212 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8215 = _T_8211 | _T_8214; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8216 = _T_8215 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8226 = _T_4732 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8227 = perr_ic_index_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8229 = _T_8227 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8230 = _T_8226 | _T_8229; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8231 = _T_8230 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8241 = _T_4733 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8242 = perr_ic_index_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8244 = _T_8242 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8245 = _T_8241 | _T_8244; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8246 = _T_8245 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8256 = _T_4734 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8257 = perr_ic_index_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8259 = _T_8257 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8260 = _T_8256 | _T_8259; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8261 = _T_8260 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8271 = _T_4735 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8272 = perr_ic_index_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8274 = _T_8272 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8275 = _T_8271 | _T_8274; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8276 = _T_8275 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8286 = _T_4736 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8287 = perr_ic_index_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8289 = _T_8287 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8290 = _T_8286 | _T_8289; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8291 = _T_8290 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8301 = _T_4737 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8302 = perr_ic_index_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8304 = _T_8302 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8305 = _T_8301 | _T_8304; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8306 = _T_8305 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8316 = _T_4738 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8317 = perr_ic_index_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8319 = _T_8317 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8320 = _T_8316 | _T_8319; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8321 = _T_8320 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8331 = _T_4739 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8332 = perr_ic_index_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8334 = _T_8332 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8335 = _T_8331 | _T_8334; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8336 = _T_8335 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8346 = _T_4740 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8347 = perr_ic_index_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8349 = _T_8347 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8350 = _T_8346 | _T_8349; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8351 = _T_8350 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8361 = _T_4741 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8362 = perr_ic_index_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8364 = _T_8362 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8365 = _T_8361 | _T_8364; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8366 = _T_8365 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8376 = _T_4742 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8377 = perr_ic_index_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8379 = _T_8377 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8380 = _T_8376 | _T_8379; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8381 = _T_8380 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8391 = _T_4743 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8392 = perr_ic_index_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8394 = _T_8392 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8395 = _T_8391 | _T_8394; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8396 = _T_8395 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8406 = _T_4744 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8407 = perr_ic_index_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8409 = _T_8407 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8410 = _T_8406 | _T_8409; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8411 = _T_8410 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8421 = _T_4745 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8422 = perr_ic_index_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8424 = _T_8422 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8425 = _T_8421 | _T_8424; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8426 = _T_8425 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8436 = _T_4746 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8437 = perr_ic_index_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8439 = _T_8437 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8440 = _T_8436 | _T_8439; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8441 = _T_8440 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8451 = _T_4747 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8452 = perr_ic_index_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 761:98]
  wire  _T_8454 = _T_8452 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8455 = _T_8451 | _T_8454; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8456 = _T_8455 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8466 = _T_4716 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8469 = _T_7987 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8470 = _T_8466 | _T_8469; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8471 = _T_8470 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8481 = _T_4717 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8484 = _T_8002 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8485 = _T_8481 | _T_8484; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8486 = _T_8485 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8496 = _T_4718 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8499 = _T_8017 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8500 = _T_8496 | _T_8499; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8501 = _T_8500 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8511 = _T_4719 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8514 = _T_8032 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8515 = _T_8511 | _T_8514; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8516 = _T_8515 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8526 = _T_4720 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8529 = _T_8047 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8530 = _T_8526 | _T_8529; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8531 = _T_8530 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8541 = _T_4721 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8544 = _T_8062 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8545 = _T_8541 | _T_8544; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8546 = _T_8545 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8556 = _T_4722 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8559 = _T_8077 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8560 = _T_8556 | _T_8559; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8561 = _T_8560 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8571 = _T_4723 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8574 = _T_8092 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8575 = _T_8571 | _T_8574; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8576 = _T_8575 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8586 = _T_4724 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8589 = _T_8107 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8590 = _T_8586 | _T_8589; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8591 = _T_8590 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8601 = _T_4725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8604 = _T_8122 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8605 = _T_8601 | _T_8604; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8606 = _T_8605 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8616 = _T_4726 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8619 = _T_8137 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8620 = _T_8616 | _T_8619; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8621 = _T_8620 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8631 = _T_4727 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8634 = _T_8152 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8635 = _T_8631 | _T_8634; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8636 = _T_8635 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8646 = _T_4728 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8649 = _T_8167 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8650 = _T_8646 | _T_8649; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8651 = _T_8650 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8661 = _T_4729 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8664 = _T_8182 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8665 = _T_8661 | _T_8664; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8666 = _T_8665 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8676 = _T_4730 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8679 = _T_8197 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8680 = _T_8676 | _T_8679; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8681 = _T_8680 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8691 = _T_4731 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8694 = _T_8212 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8695 = _T_8691 | _T_8694; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8696 = _T_8695 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8706 = _T_4732 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8709 = _T_8227 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8710 = _T_8706 | _T_8709; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8711 = _T_8710 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8721 = _T_4733 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8724 = _T_8242 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8725 = _T_8721 | _T_8724; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8726 = _T_8725 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8736 = _T_4734 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8739 = _T_8257 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8740 = _T_8736 | _T_8739; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8741 = _T_8740 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8751 = _T_4735 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8754 = _T_8272 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8755 = _T_8751 | _T_8754; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8756 = _T_8755 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8766 = _T_4736 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8769 = _T_8287 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8770 = _T_8766 | _T_8769; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8771 = _T_8770 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8781 = _T_4737 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8784 = _T_8302 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8785 = _T_8781 | _T_8784; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8786 = _T_8785 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8796 = _T_4738 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8799 = _T_8317 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8800 = _T_8796 | _T_8799; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8801 = _T_8800 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8811 = _T_4739 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8814 = _T_8332 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8815 = _T_8811 | _T_8814; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8816 = _T_8815 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8826 = _T_4740 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8829 = _T_8347 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8830 = _T_8826 | _T_8829; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8831 = _T_8830 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8841 = _T_4741 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8844 = _T_8362 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8845 = _T_8841 | _T_8844; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8846 = _T_8845 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8856 = _T_4742 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8859 = _T_8377 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8860 = _T_8856 | _T_8859; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8861 = _T_8860 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8871 = _T_4743 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8874 = _T_8392 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8875 = _T_8871 | _T_8874; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8876 = _T_8875 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8886 = _T_4744 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8889 = _T_8407 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8890 = _T_8886 | _T_8889; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8891 = _T_8890 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8901 = _T_4745 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8904 = _T_8422 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8905 = _T_8901 | _T_8904; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8906 = _T_8905 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8916 = _T_4746 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8919 = _T_8437 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8920 = _T_8916 | _T_8919; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8921 = _T_8920 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_8931 = _T_4747 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:55]
  wire  _T_8934 = _T_8452 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:120]
  wire  _T_8935 = _T_8931 | _T_8934; // @[el2_ifu_mem_ctl.scala 761:77]
  wire  _T_8936 = _T_8935 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:143]
  wire  _T_9738 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 816:63]
  wire  _T_9739 = _T_9738 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 816:85]
  wire [1:0] _T_9741 = _T_9739 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9748; // @[el2_ifu_mem_ctl.scala 821:57]
  reg  _T_9749; // @[el2_ifu_mem_ctl.scala 822:56]
  reg  _T_9750; // @[el2_ifu_mem_ctl.scala 823:59]
  wire  _T_9751 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 824:80]
  wire  _T_9752 = ifu_bus_arvalid_ff & _T_9751; // @[el2_ifu_mem_ctl.scala 824:78]
  reg  _T_9754; // @[el2_ifu_mem_ctl.scala 824:58]
  reg  _T_9755; // @[el2_ifu_mem_ctl.scala 825:58]
  wire  _T_9758 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 832:71]
  wire  _T_9760 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 832:124]
  wire  _T_9762 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 833:50]
  wire  _T_9764 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 833:103]
  wire [3:0] _T_9767 = {_T_9758,_T_9760,_T_9762,_T_9764}; // @[Cat.scala 29:58]
  reg  _T_9776; // @[Reg.scala 27:20]
  wire [31:0] _T_9786 = {io_ifc_fetch_addr_bf,1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_9787 = _T_9786 | 32'h7fffffff; // @[el2_ifu_mem_ctl.scala 841:63]
  wire  _T_9789 = _T_9787 == 32'h7fffffff; // @[el2_ifu_mem_ctl.scala 841:94]
  wire [31:0] _T_9793 = _T_9786 | 32'h3fffffff; // @[el2_ifu_mem_ctl.scala 842:63]
  wire  _T_9795 = _T_9793 == 32'hffffffff; // @[el2_ifu_mem_ctl.scala 842:94]
  wire  _T_9797 = _T_9789 | _T_9795; // @[el2_ifu_mem_ctl.scala 841:160]
  wire [31:0] _T_9799 = _T_9786 | 32'h1fffffff; // @[el2_ifu_mem_ctl.scala 843:63]
  wire  _T_9801 = _T_9799 == 32'hbfffffff; // @[el2_ifu_mem_ctl.scala 843:94]
  wire  _T_9803 = _T_9797 | _T_9801; // @[el2_ifu_mem_ctl.scala 842:160]
  wire [31:0] _T_9805 = _T_9786 | 32'hfffffff; // @[el2_ifu_mem_ctl.scala 844:63]
  wire  _T_9807 = _T_9805 == 32'h8fffffff; // @[el2_ifu_mem_ctl.scala 844:94]
  wire  ifc_region_acc_okay = _T_9803 | _T_9807; // @[el2_ifu_mem_ctl.scala 843:160]
  wire  _T_9834 = ~ifc_region_acc_okay; // @[el2_ifu_mem_ctl.scala 849:65]
  wire  _T_9835 = _T_3888 & _T_9834; // @[el2_ifu_mem_ctl.scala 849:63]
  wire  ifc_region_acc_fault_memory_bf = _T_9835 & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 849:86]
  rvclkhdr rvclkhdr ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  rvclkhdr rvclkhdr_26 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_26_io_l1clk),
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en),
    .io_scan_mode(rvclkhdr_26_io_scan_mode)
  );
  rvclkhdr rvclkhdr_27 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_27_io_l1clk),
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en),
    .io_scan_mode(rvclkhdr_27_io_scan_mode)
  );
  rvclkhdr rvclkhdr_28 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_28_io_l1clk),
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en),
    .io_scan_mode(rvclkhdr_28_io_scan_mode)
  );
  rvclkhdr rvclkhdr_29 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_29_io_l1clk),
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en),
    .io_scan_mode(rvclkhdr_29_io_scan_mode)
  );
  rvclkhdr rvclkhdr_30 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_30_io_l1clk),
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en),
    .io_scan_mode(rvclkhdr_30_io_scan_mode)
  );
  rvclkhdr rvclkhdr_31 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_31_io_l1clk),
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en),
    .io_scan_mode(rvclkhdr_31_io_scan_mode)
  );
  rvclkhdr rvclkhdr_32 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_32_io_l1clk),
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en),
    .io_scan_mode(rvclkhdr_32_io_scan_mode)
  );
  rvclkhdr rvclkhdr_33 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_33_io_l1clk),
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en),
    .io_scan_mode(rvclkhdr_33_io_scan_mode)
  );
  rvclkhdr rvclkhdr_34 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_34_io_l1clk),
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en),
    .io_scan_mode(rvclkhdr_34_io_scan_mode)
  );
  rvclkhdr rvclkhdr_35 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_35_io_l1clk),
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en),
    .io_scan_mode(rvclkhdr_35_io_scan_mode)
  );
  rvclkhdr rvclkhdr_36 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_36_io_l1clk),
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en),
    .io_scan_mode(rvclkhdr_36_io_scan_mode)
  );
  rvclkhdr rvclkhdr_37 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_37_io_l1clk),
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en),
    .io_scan_mode(rvclkhdr_37_io_scan_mode)
  );
  rvclkhdr rvclkhdr_38 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_38_io_l1clk),
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en),
    .io_scan_mode(rvclkhdr_38_io_scan_mode)
  );
  rvclkhdr rvclkhdr_39 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_39_io_l1clk),
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en),
    .io_scan_mode(rvclkhdr_39_io_scan_mode)
  );
  rvclkhdr rvclkhdr_40 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_40_io_l1clk),
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en),
    .io_scan_mode(rvclkhdr_40_io_scan_mode)
  );
  rvclkhdr rvclkhdr_41 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_41_io_l1clk),
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en),
    .io_scan_mode(rvclkhdr_41_io_scan_mode)
  );
  rvclkhdr rvclkhdr_42 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_42_io_l1clk),
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en),
    .io_scan_mode(rvclkhdr_42_io_scan_mode)
  );
  rvclkhdr rvclkhdr_43 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_43_io_l1clk),
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en),
    .io_scan_mode(rvclkhdr_43_io_scan_mode)
  );
  rvclkhdr rvclkhdr_44 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_44_io_l1clk),
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en),
    .io_scan_mode(rvclkhdr_44_io_scan_mode)
  );
  rvclkhdr rvclkhdr_45 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_45_io_l1clk),
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en),
    .io_scan_mode(rvclkhdr_45_io_scan_mode)
  );
  rvclkhdr rvclkhdr_46 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_46_io_l1clk),
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en),
    .io_scan_mode(rvclkhdr_46_io_scan_mode)
  );
  rvclkhdr rvclkhdr_47 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_47_io_l1clk),
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en),
    .io_scan_mode(rvclkhdr_47_io_scan_mode)
  );
  rvclkhdr rvclkhdr_48 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_48_io_l1clk),
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en),
    .io_scan_mode(rvclkhdr_48_io_scan_mode)
  );
  rvclkhdr rvclkhdr_49 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_49_io_l1clk),
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en),
    .io_scan_mode(rvclkhdr_49_io_scan_mode)
  );
  rvclkhdr rvclkhdr_50 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_50_io_l1clk),
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en),
    .io_scan_mode(rvclkhdr_50_io_scan_mode)
  );
  rvclkhdr rvclkhdr_51 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_51_io_l1clk),
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en),
    .io_scan_mode(rvclkhdr_51_io_scan_mode)
  );
  rvclkhdr rvclkhdr_52 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_52_io_l1clk),
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en),
    .io_scan_mode(rvclkhdr_52_io_scan_mode)
  );
  rvclkhdr rvclkhdr_53 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_53_io_l1clk),
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en),
    .io_scan_mode(rvclkhdr_53_io_scan_mode)
  );
  rvclkhdr rvclkhdr_54 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_54_io_l1clk),
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en),
    .io_scan_mode(rvclkhdr_54_io_scan_mode)
  );
  rvclkhdr rvclkhdr_55 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_55_io_l1clk),
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en),
    .io_scan_mode(rvclkhdr_55_io_scan_mode)
  );
  rvclkhdr rvclkhdr_56 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_56_io_l1clk),
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en),
    .io_scan_mode(rvclkhdr_56_io_scan_mode)
  );
  rvclkhdr rvclkhdr_57 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_57_io_l1clk),
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en),
    .io_scan_mode(rvclkhdr_57_io_scan_mode)
  );
  rvclkhdr rvclkhdr_58 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_58_io_l1clk),
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en),
    .io_scan_mode(rvclkhdr_58_io_scan_mode)
  );
  rvclkhdr rvclkhdr_59 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_59_io_l1clk),
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en),
    .io_scan_mode(rvclkhdr_59_io_scan_mode)
  );
  rvclkhdr rvclkhdr_60 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_60_io_l1clk),
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en),
    .io_scan_mode(rvclkhdr_60_io_scan_mode)
  );
  rvclkhdr rvclkhdr_61 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_61_io_l1clk),
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en),
    .io_scan_mode(rvclkhdr_61_io_scan_mode)
  );
  rvclkhdr rvclkhdr_62 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_62_io_l1clk),
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en),
    .io_scan_mode(rvclkhdr_62_io_scan_mode)
  );
  rvclkhdr rvclkhdr_63 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_63_io_l1clk),
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en),
    .io_scan_mode(rvclkhdr_63_io_scan_mode)
  );
  rvclkhdr rvclkhdr_64 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_64_io_l1clk),
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en),
    .io_scan_mode(rvclkhdr_64_io_scan_mode)
  );
  rvclkhdr rvclkhdr_65 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_65_io_l1clk),
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en),
    .io_scan_mode(rvclkhdr_65_io_scan_mode)
  );
  rvclkhdr rvclkhdr_66 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_66_io_l1clk),
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en),
    .io_scan_mode(rvclkhdr_66_io_scan_mode)
  );
  rvclkhdr rvclkhdr_67 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_67_io_l1clk),
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en),
    .io_scan_mode(rvclkhdr_67_io_scan_mode)
  );
  rvclkhdr rvclkhdr_68 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_68_io_l1clk),
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en),
    .io_scan_mode(rvclkhdr_68_io_scan_mode)
  );
  rvclkhdr rvclkhdr_69 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_69_io_l1clk),
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en),
    .io_scan_mode(rvclkhdr_69_io_scan_mode)
  );
  rvclkhdr rvclkhdr_70 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_70_io_l1clk),
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en),
    .io_scan_mode(rvclkhdr_70_io_scan_mode)
  );
  rvclkhdr rvclkhdr_71 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_71_io_l1clk),
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en),
    .io_scan_mode(rvclkhdr_71_io_scan_mode)
  );
  rvclkhdr rvclkhdr_72 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_72_io_l1clk),
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en),
    .io_scan_mode(rvclkhdr_72_io_scan_mode)
  );
  rvclkhdr rvclkhdr_73 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_73_io_l1clk),
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en),
    .io_scan_mode(rvclkhdr_73_io_scan_mode)
  );
  rvclkhdr rvclkhdr_74 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_74_io_l1clk),
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en),
    .io_scan_mode(rvclkhdr_74_io_scan_mode)
  );
  rvclkhdr rvclkhdr_75 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_75_io_l1clk),
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en),
    .io_scan_mode(rvclkhdr_75_io_scan_mode)
  );
  rvclkhdr rvclkhdr_76 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_76_io_l1clk),
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en),
    .io_scan_mode(rvclkhdr_76_io_scan_mode)
  );
  rvclkhdr rvclkhdr_77 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_77_io_l1clk),
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en),
    .io_scan_mode(rvclkhdr_77_io_scan_mode)
  );
  rvclkhdr rvclkhdr_78 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_78_io_l1clk),
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en),
    .io_scan_mode(rvclkhdr_78_io_scan_mode)
  );
  rvclkhdr rvclkhdr_79 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_79_io_l1clk),
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en),
    .io_scan_mode(rvclkhdr_79_io_scan_mode)
  );
  rvclkhdr rvclkhdr_80 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_80_io_l1clk),
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en),
    .io_scan_mode(rvclkhdr_80_io_scan_mode)
  );
  rvclkhdr rvclkhdr_81 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_81_io_l1clk),
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en),
    .io_scan_mode(rvclkhdr_81_io_scan_mode)
  );
  rvclkhdr rvclkhdr_82 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_82_io_l1clk),
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en),
    .io_scan_mode(rvclkhdr_82_io_scan_mode)
  );
  rvclkhdr rvclkhdr_83 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_83_io_l1clk),
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en),
    .io_scan_mode(rvclkhdr_83_io_scan_mode)
  );
  rvclkhdr rvclkhdr_84 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_84_io_l1clk),
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en),
    .io_scan_mode(rvclkhdr_84_io_scan_mode)
  );
  rvclkhdr rvclkhdr_85 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_85_io_l1clk),
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en),
    .io_scan_mode(rvclkhdr_85_io_scan_mode)
  );
  rvclkhdr rvclkhdr_86 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_86_io_l1clk),
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en),
    .io_scan_mode(rvclkhdr_86_io_scan_mode)
  );
  rvclkhdr rvclkhdr_87 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_87_io_l1clk),
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en),
    .io_scan_mode(rvclkhdr_87_io_scan_mode)
  );
  rvclkhdr rvclkhdr_88 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_88_io_l1clk),
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en),
    .io_scan_mode(rvclkhdr_88_io_scan_mode)
  );
  rvclkhdr rvclkhdr_89 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_89_io_l1clk),
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en),
    .io_scan_mode(rvclkhdr_89_io_scan_mode)
  );
  rvclkhdr rvclkhdr_90 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_90_io_l1clk),
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en),
    .io_scan_mode(rvclkhdr_90_io_scan_mode)
  );
  rvclkhdr rvclkhdr_91 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_91_io_l1clk),
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en),
    .io_scan_mode(rvclkhdr_91_io_scan_mode)
  );
  rvclkhdr rvclkhdr_92 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_92_io_l1clk),
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en),
    .io_scan_mode(rvclkhdr_92_io_scan_mode)
  );
  rvclkhdr rvclkhdr_93 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_93_io_l1clk),
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en),
    .io_scan_mode(rvclkhdr_93_io_scan_mode)
  );
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 330:26]
  assign io_ifu_ic_mb_empty = _T_328 | _T_231; // @[el2_ifu_mem_ctl.scala 329:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 193:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3937; // @[el2_ifu_mem_ctl.scala 704:21]
  assign io_ifu_pmu_ic_miss = _T_9748; // @[el2_ifu_mem_ctl.scala 821:22]
  assign io_ifu_pmu_ic_hit = _T_9749; // @[el2_ifu_mem_ctl.scala 822:21]
  assign io_ifu_pmu_bus_error = _T_9750; // @[el2_ifu_mem_ctl.scala 823:24]
  assign io_ifu_pmu_bus_busy = _T_9754; // @[el2_ifu_mem_ctl.scala 824:23]
  assign io_ifu_pmu_bus_trxn = _T_9755; // @[el2_ifu_mem_ctl.scala 825:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 144:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 143:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 138:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 142:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 140:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 151:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 153:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 148:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 146:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 139:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 137:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 135:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 136:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 145:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 154:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 149:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 565:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2559; // @[el2_ifu_mem_ctl.scala 566:19]
  assign io_ifu_axi_araddr = _T_2561 & _T_2563; // @[el2_ifu_mem_ctl.scala 567:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 570:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 150:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 568:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 571:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 141:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 569:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 152:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 147:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 572:21]
  assign io_iccm_dma_ecc_error = iccm_dma_ecc_error; // @[el2_ifu_mem_ctl.scala 663:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 661:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 665:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 656:20]
  assign io_iccm_ready = _T_2657 & _T_2651; // @[el2_ifu_mem_ctl.scala 635:17]
  assign io_ic_rw_addr = _T_340 | _T_341; // @[el2_ifu_mem_ctl.scala 339:17]
  assign io_ic_wr_en = bus_ic_wr_en & _T_3923; // @[el2_ifu_mem_ctl.scala 703:15]
  assign io_ic_rd_en = _T_3915 | _T_3920; // @[el2_ifu_mem_ctl.scala 694:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 346:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 346:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 347:23]
  assign io_ifu_ic_debug_rd_data = _T_1211; // @[el2_ifu_mem_ctl.scala 355:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 828:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 830:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 831:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 829:25]
  assign io_ic_debug_way = _T_9767[1:0]; // @[el2_ifu_mem_ctl.scala 832:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9741; // @[el2_ifu_mem_ctl.scala 816:19]
  assign io_iccm_rw_addr = _T_3061 ? io_dma_mem_addr[15:1] : _T_3068; // @[el2_ifu_mem_ctl.scala 667:19]
  assign io_iccm_wren = _T_2661 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 637:16]
  assign io_iccm_rden = _T_2665 | _T_2666; // @[el2_ifu_mem_ctl.scala 638:16]
  assign io_iccm_wr_data = _T_3043 ? _T_3044 : _T_3051; // @[el2_ifu_mem_ctl.scala 644:19]
  assign io_iccm_wr_size = _T_2671 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 640:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 290:15]
  assign io_ic_access_fault_f = _T_2443 & _T_319; // @[el2_ifu_mem_ctl.scala 387:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1273; // @[el2_ifu_mem_ctl.scala 388:29]
  assign io_iccm_rd_ecc_single_err = _T_3860 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 680:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 681:29]
  assign io_ic_error_start = _T_1199 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 349:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 192:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 191:24]
  assign io_ic_fetch_val_f = {_T_1281,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 391:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 384:16]
  assign io_ic_premux_data = ic_premux_data_temp[63:0]; // @[el2_ifu_mem_ctl.scala 381:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 382:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_9776; // @[el2_ifu_mem_ctl.scala 839:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2448; // @[el2_ifu_mem_ctl.scala 482:27]
  assign io_iccm_correction_state = _T_2477 ? 1'h0 : _GEN_43; // @[el2_ifu_mem_ctl.scala 517:28 el2_ifu_mem_ctl.scala 530:32 el2_ifu_mem_ctl.scala 537:32 el2_ifu_mem_ctl.scala 544:32]
  assign rvclkhdr_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_io_en = ic_debug_rd_en_ff; // @[el2_lib.scala 485:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_1_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_1_io_en = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_lib.scala 485:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_2_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_2_io_en = _T_2 | scnd_miss_req; // @[el2_lib.scala 485:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_3_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_3_io_en = _T_309 | io_dec_tlu_force_halt; // @[el2_lib.scala 485:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_4_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_4_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_5_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_5_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_6_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_6_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_7_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_7_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_8_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_8_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_9_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_9_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_10_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_10_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_11_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_11_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_12_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_12_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_13_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_13_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_14_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_14_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_15_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_15_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_16_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_16_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_17_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_17_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_18_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_18_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_19_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_19_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_20_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_20_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_21_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_21_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_22_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_22_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_23_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_23_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_24_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_24_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_25_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_25_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_26_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_26_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_26_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_27_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_27_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_27_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_28_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_28_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_28_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_29_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_29_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_29_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_30_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_30_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_30_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_31_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_31_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_31_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_32_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_32_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_32_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_33_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_33_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_33_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_34_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_34_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_34_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_35_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_35_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_35_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_36_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_36_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_36_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_37_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_37_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_37_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_38_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_38_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_38_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_39_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_39_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_39_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_40_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_40_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_40_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_41_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_41_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_41_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_42_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_42_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_42_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_43_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_43_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_43_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_44_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_44_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_44_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_45_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_45_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_45_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_46_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_46_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_46_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_47_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_47_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_47_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_48_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_48_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_48_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_49_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_49_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_49_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_50_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_50_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_50_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_51_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_51_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_51_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_52_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_52_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_52_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_53_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_53_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_53_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_54_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_54_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_54_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_55_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_55_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_55_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_56_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_56_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_56_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_57_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_57_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_57_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_58_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_58_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_58_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_59_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_59_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_59_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_60_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_60_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_60_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_61_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_61_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_61_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_62_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_62_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_62_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_63_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_63_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_63_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_64_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_64_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_64_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_65_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_65_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_65_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_66_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_66_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_66_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_67_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_67_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_67_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_68_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_68_io_en = io_ifu_bus_clk_en; // @[el2_lib.scala 485:16]
  assign rvclkhdr_68_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_69_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_69_io_en = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_lib.scala 485:16]
  assign rvclkhdr_69_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_70_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_70_io_en = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_lib.scala 485:16]
  assign rvclkhdr_70_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_71_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_71_io_en = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_lib.scala 485:16]
  assign rvclkhdr_71_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_72_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_72_io_en = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_lib.scala 485:16]
  assign rvclkhdr_72_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_73_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_73_io_en = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_lib.scala 485:16]
  assign rvclkhdr_73_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_74_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_74_io_en = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_lib.scala 485:16]
  assign rvclkhdr_74_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_75_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_75_io_en = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_lib.scala 485:16]
  assign rvclkhdr_75_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_76_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_76_io_en = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_lib.scala 485:16]
  assign rvclkhdr_76_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_77_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_77_io_en = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_lib.scala 485:16]
  assign rvclkhdr_77_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_78_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_78_io_en = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_lib.scala 485:16]
  assign rvclkhdr_78_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_79_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_79_io_en = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_lib.scala 485:16]
  assign rvclkhdr_79_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_80_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_80_io_en = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_lib.scala 485:16]
  assign rvclkhdr_80_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_81_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_81_io_en = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_lib.scala 485:16]
  assign rvclkhdr_81_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_82_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_82_io_en = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_lib.scala 485:16]
  assign rvclkhdr_82_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_83_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_83_io_en = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_lib.scala 485:16]
  assign rvclkhdr_83_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_84_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_84_io_en = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_lib.scala 485:16]
  assign rvclkhdr_84_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_85_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_85_io_en = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_lib.scala 485:16]
  assign rvclkhdr_85_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_86_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_86_io_en = tag_valid_clken_0[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_86_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_87_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_87_io_en = tag_valid_clken_0[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_87_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_88_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_88_io_en = tag_valid_clken_1[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_88_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_89_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_89_io_en = tag_valid_clken_1[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_89_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_90_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_90_io_en = tag_valid_clken_2[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_90_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_91_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_91_io_en = tag_valid_clken_2[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_91_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_92_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_92_io_en = tag_valid_clken_3[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_92_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_93_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_93_io_en = tag_valid_clken_3[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_93_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_11 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_17 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_18 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_19 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_20 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_21 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_23 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_24 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_25 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_26 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_27 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_29 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_30 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_32 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_33 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_34 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_35 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_36 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_37 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_38 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_39 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_40 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_41 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_42 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_43 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_44 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_45 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_46 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_47 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_48 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_49 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_50 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_51 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_52 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_53 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_54 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_55 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_56 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_57 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_58 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_59 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_60 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_61 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_62 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_63 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_64 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_65 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_66 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_67 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_68 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_69 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_70 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_71 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_72 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_73 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_74 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_75 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_76 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_77 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_78 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_79 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_80 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_81 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_82 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_83 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_84 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_85 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_86 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_87 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_88 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_89 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_90 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_91 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_92 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_93 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_94 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_95 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_96 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_97 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_98 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_99 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_100 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_101 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_102 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_103 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_104 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_105 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_106 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_107 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_108 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_109 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_110 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_111 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_112 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_113 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_114 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_115 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_116 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_117 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_118 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_119 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_120 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_121 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_out_122 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way_status_out_123 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way_status_out_124 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way_status_out_125 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way_status_out_126 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way_status_out_127 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagv_mb_scnd_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_152[30:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  reset_ic_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  miss_addr = _RAND_160[25:0];
  _RAND_161 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_441[0:0];
  _RAND_442 = {3{`RANDOM}};
  _T_1211 = _RAND_442[70:0];
  _RAND_443 = {1{`RANDOM}};
  ifc_region_acc_fault_memory_f = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_444[6:0];
  _RAND_445 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  bus_cmd_req_hold = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_448[2:0];
  _RAND_449 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_451[0:0];
  _RAND_452 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_452[38:0];
  _RAND_453 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_454[2:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_dma_rtag_temp = _RAND_455[2:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_dma_rvalid_temp = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_dma_ecc_error = _RAND_457[0:0];
  _RAND_458 = {2{`RANDOM}};
  iccm_dma_rdata_temp = _RAND_458[63:0];
  _RAND_459 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_459[13:0];
  _RAND_460 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_461[13:0];
  _RAND_462 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_462[6:0];
  _RAND_463 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  way_status_new_ff = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  ic_valid_ff = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_9748 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_9749 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_9750 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  _T_9754 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  _T_9755 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  _T_9776 = _RAND_472[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    flush_final_f = 1'h0;
  end
  if (reset) begin
    ifc_fetch_req_f_raw = 1'h0;
  end
  if (reset) begin
    miss_state = 3'h0;
  end
  if (reset) begin
    scnd_miss_req_q = 1'h0;
  end
  if (reset) begin
    ifu_fetch_addr_int_f = 31'h0;
  end
  if (reset) begin
    ifc_iccm_access_f = 1'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_in = 1'h0;
  end
  if (reset) begin
    dma_iccm_req_f = 1'h0;
  end
  if (reset) begin
    perr_state = 3'h0;
  end
  if (reset) begin
    err_stop_state = 2'h0;
  end
  if (reset) begin
    reset_all_tags = 1'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_final_f = 1'h0;
  end
  if (reset) begin
    ifu_bus_rvalid_unq_ff = 1'h0;
  end
  if (reset) begin
    bus_ifu_bus_clk_en_ff = 1'h0;
  end
  if (reset) begin
    uncacheable_miss_ff = 1'h0;
  end
  if (reset) begin
    bus_data_beat_count = 3'h0;
  end
  if (reset) begin
    ic_miss_buff_data_valid = 8'h0;
  end
  if (reset) begin
    last_data_recieved_ff = 1'h0;
  end
  if (reset) begin
    sel_mb_addr_ff = 1'h0;
  end
  if (reset) begin
    way_status_mb_scnd_ff = 1'h0;
  end
  if (reset) begin
    ifu_ic_rw_int_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_out_0 = 1'h0;
  end
  if (reset) begin
    way_status_out_1 = 1'h0;
  end
  if (reset) begin
    way_status_out_2 = 1'h0;
  end
  if (reset) begin
    way_status_out_3 = 1'h0;
  end
  if (reset) begin
    way_status_out_4 = 1'h0;
  end
  if (reset) begin
    way_status_out_5 = 1'h0;
  end
  if (reset) begin
    way_status_out_6 = 1'h0;
  end
  if (reset) begin
    way_status_out_7 = 1'h0;
  end
  if (reset) begin
    way_status_out_8 = 1'h0;
  end
  if (reset) begin
    way_status_out_9 = 1'h0;
  end
  if (reset) begin
    way_status_out_10 = 1'h0;
  end
  if (reset) begin
    way_status_out_11 = 1'h0;
  end
  if (reset) begin
    way_status_out_12 = 1'h0;
  end
  if (reset) begin
    way_status_out_13 = 1'h0;
  end
  if (reset) begin
    way_status_out_14 = 1'h0;
  end
  if (reset) begin
    way_status_out_15 = 1'h0;
  end
  if (reset) begin
    way_status_out_16 = 1'h0;
  end
  if (reset) begin
    way_status_out_17 = 1'h0;
  end
  if (reset) begin
    way_status_out_18 = 1'h0;
  end
  if (reset) begin
    way_status_out_19 = 1'h0;
  end
  if (reset) begin
    way_status_out_20 = 1'h0;
  end
  if (reset) begin
    way_status_out_21 = 1'h0;
  end
  if (reset) begin
    way_status_out_22 = 1'h0;
  end
  if (reset) begin
    way_status_out_23 = 1'h0;
  end
  if (reset) begin
    way_status_out_24 = 1'h0;
  end
  if (reset) begin
    way_status_out_25 = 1'h0;
  end
  if (reset) begin
    way_status_out_26 = 1'h0;
  end
  if (reset) begin
    way_status_out_27 = 1'h0;
  end
  if (reset) begin
    way_status_out_28 = 1'h0;
  end
  if (reset) begin
    way_status_out_29 = 1'h0;
  end
  if (reset) begin
    way_status_out_30 = 1'h0;
  end
  if (reset) begin
    way_status_out_31 = 1'h0;
  end
  if (reset) begin
    way_status_out_32 = 1'h0;
  end
  if (reset) begin
    way_status_out_33 = 1'h0;
  end
  if (reset) begin
    way_status_out_34 = 1'h0;
  end
  if (reset) begin
    way_status_out_35 = 1'h0;
  end
  if (reset) begin
    way_status_out_36 = 1'h0;
  end
  if (reset) begin
    way_status_out_37 = 1'h0;
  end
  if (reset) begin
    way_status_out_38 = 1'h0;
  end
  if (reset) begin
    way_status_out_39 = 1'h0;
  end
  if (reset) begin
    way_status_out_40 = 1'h0;
  end
  if (reset) begin
    way_status_out_41 = 1'h0;
  end
  if (reset) begin
    way_status_out_42 = 1'h0;
  end
  if (reset) begin
    way_status_out_43 = 1'h0;
  end
  if (reset) begin
    way_status_out_44 = 1'h0;
  end
  if (reset) begin
    way_status_out_45 = 1'h0;
  end
  if (reset) begin
    way_status_out_46 = 1'h0;
  end
  if (reset) begin
    way_status_out_47 = 1'h0;
  end
  if (reset) begin
    way_status_out_48 = 1'h0;
  end
  if (reset) begin
    way_status_out_49 = 1'h0;
  end
  if (reset) begin
    way_status_out_50 = 1'h0;
  end
  if (reset) begin
    way_status_out_51 = 1'h0;
  end
  if (reset) begin
    way_status_out_52 = 1'h0;
  end
  if (reset) begin
    way_status_out_53 = 1'h0;
  end
  if (reset) begin
    way_status_out_54 = 1'h0;
  end
  if (reset) begin
    way_status_out_55 = 1'h0;
  end
  if (reset) begin
    way_status_out_56 = 1'h0;
  end
  if (reset) begin
    way_status_out_57 = 1'h0;
  end
  if (reset) begin
    way_status_out_58 = 1'h0;
  end
  if (reset) begin
    way_status_out_59 = 1'h0;
  end
  if (reset) begin
    way_status_out_60 = 1'h0;
  end
  if (reset) begin
    way_status_out_61 = 1'h0;
  end
  if (reset) begin
    way_status_out_62 = 1'h0;
  end
  if (reset) begin
    way_status_out_63 = 1'h0;
  end
  if (reset) begin
    way_status_out_64 = 1'h0;
  end
  if (reset) begin
    way_status_out_65 = 1'h0;
  end
  if (reset) begin
    way_status_out_66 = 1'h0;
  end
  if (reset) begin
    way_status_out_67 = 1'h0;
  end
  if (reset) begin
    way_status_out_68 = 1'h0;
  end
  if (reset) begin
    way_status_out_69 = 1'h0;
  end
  if (reset) begin
    way_status_out_70 = 1'h0;
  end
  if (reset) begin
    way_status_out_71 = 1'h0;
  end
  if (reset) begin
    way_status_out_72 = 1'h0;
  end
  if (reset) begin
    way_status_out_73 = 1'h0;
  end
  if (reset) begin
    way_status_out_74 = 1'h0;
  end
  if (reset) begin
    way_status_out_75 = 1'h0;
  end
  if (reset) begin
    way_status_out_76 = 1'h0;
  end
  if (reset) begin
    way_status_out_77 = 1'h0;
  end
  if (reset) begin
    way_status_out_78 = 1'h0;
  end
  if (reset) begin
    way_status_out_79 = 1'h0;
  end
  if (reset) begin
    way_status_out_80 = 1'h0;
  end
  if (reset) begin
    way_status_out_81 = 1'h0;
  end
  if (reset) begin
    way_status_out_82 = 1'h0;
  end
  if (reset) begin
    way_status_out_83 = 1'h0;
  end
  if (reset) begin
    way_status_out_84 = 1'h0;
  end
  if (reset) begin
    way_status_out_85 = 1'h0;
  end
  if (reset) begin
    way_status_out_86 = 1'h0;
  end
  if (reset) begin
    way_status_out_87 = 1'h0;
  end
  if (reset) begin
    way_status_out_88 = 1'h0;
  end
  if (reset) begin
    way_status_out_89 = 1'h0;
  end
  if (reset) begin
    way_status_out_90 = 1'h0;
  end
  if (reset) begin
    way_status_out_91 = 1'h0;
  end
  if (reset) begin
    way_status_out_92 = 1'h0;
  end
  if (reset) begin
    way_status_out_93 = 1'h0;
  end
  if (reset) begin
    way_status_out_94 = 1'h0;
  end
  if (reset) begin
    way_status_out_95 = 1'h0;
  end
  if (reset) begin
    way_status_out_96 = 1'h0;
  end
  if (reset) begin
    way_status_out_97 = 1'h0;
  end
  if (reset) begin
    way_status_out_98 = 1'h0;
  end
  if (reset) begin
    way_status_out_99 = 1'h0;
  end
  if (reset) begin
    way_status_out_100 = 1'h0;
  end
  if (reset) begin
    way_status_out_101 = 1'h0;
  end
  if (reset) begin
    way_status_out_102 = 1'h0;
  end
  if (reset) begin
    way_status_out_103 = 1'h0;
  end
  if (reset) begin
    way_status_out_104 = 1'h0;
  end
  if (reset) begin
    way_status_out_105 = 1'h0;
  end
  if (reset) begin
    way_status_out_106 = 1'h0;
  end
  if (reset) begin
    way_status_out_107 = 1'h0;
  end
  if (reset) begin
    way_status_out_108 = 1'h0;
  end
  if (reset) begin
    way_status_out_109 = 1'h0;
  end
  if (reset) begin
    way_status_out_110 = 1'h0;
  end
  if (reset) begin
    way_status_out_111 = 1'h0;
  end
  if (reset) begin
    way_status_out_112 = 1'h0;
  end
  if (reset) begin
    way_status_out_113 = 1'h0;
  end
  if (reset) begin
    way_status_out_114 = 1'h0;
  end
  if (reset) begin
    way_status_out_115 = 1'h0;
  end
  if (reset) begin
    way_status_out_116 = 1'h0;
  end
  if (reset) begin
    way_status_out_117 = 1'h0;
  end
  if (reset) begin
    way_status_out_118 = 1'h0;
  end
  if (reset) begin
    way_status_out_119 = 1'h0;
  end
  if (reset) begin
    way_status_out_120 = 1'h0;
  end
  if (reset) begin
    way_status_out_121 = 1'h0;
  end
  if (reset) begin
    way_status_out_122 = 1'h0;
  end
  if (reset) begin
    way_status_out_123 = 1'h0;
  end
  if (reset) begin
    way_status_out_124 = 1'h0;
  end
  if (reset) begin
    way_status_out_125 = 1'h0;
  end
  if (reset) begin
    way_status_out_126 = 1'h0;
  end
  if (reset) begin
    way_status_out_127 = 1'h0;
  end
  if (reset) begin
    tagv_mb_scnd_ff = 2'h0;
  end
  if (reset) begin
    uncacheable_miss_scnd_ff = 1'h0;
  end
  if (reset) begin
    imb_scnd_ff = 31'h0;
  end
  if (reset) begin
    ifu_bus_rid_ff = 3'h0;
  end
  if (reset) begin
    ifu_bus_rresp_ff = 2'h0;
  end
  if (reset) begin
    ifu_wr_data_comb_err_ff = 1'h0;
  end
  if (reset) begin
    way_status_mb_ff = 1'h0;
  end
  if (reset) begin
    tagv_mb_ff = 2'h0;
  end
  if (reset) begin
    fetch_uncacheable_ff = 1'h0;
  end
  if (reset) begin
    miss_addr = 26'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_f = 1'h0;
  end
  if (reset) begin
    bus_rd_addr_count = 3'h0;
  end
  if (reset) begin
    ic_act_miss_f_delayed = 1'h0;
  end
  if (reset) begin
    ifu_bus_rdata_ff = 64'h0;
  end
  if (reset) begin
    ic_miss_buff_data_0 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_1 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_2 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_3 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_4 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_5 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_6 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_7 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_8 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_9 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_10 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_11 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_12 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_13 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_14 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_15 = 32'h0;
  end
  if (reset) begin
    ic_crit_wd_rdy_new_ff = 1'h0;
  end
  if (reset) begin
    ic_miss_buff_data_error = 8'h0;
  end
  if (reset) begin
    ic_debug_ict_array_sel_ff = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_127 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_127 = 1'h0;
  end
  if (reset) begin
    ic_debug_way_ff = 2'h0;
  end
  if (reset) begin
    ic_debug_rd_en_ff = 1'h0;
  end
  if (reset) begin
    _T_1211 = 71'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_memory_f = 1'h0;
  end
  if (reset) begin
    perr_ic_index_ff = 7'h0;
  end
  if (reset) begin
    dma_sb_err_state_ff = 1'h0;
  end
  if (reset) begin
    bus_cmd_req_hold = 1'h0;
  end
  if (reset) begin
    ifu_bus_cmd_valid = 1'h0;
  end
  if (reset) begin
    bus_cmd_beat_count = 3'h0;
  end
  if (reset) begin
    ifu_bus_arready_unq_ff = 1'h0;
  end
  if (reset) begin
    ifu_bus_arvalid_ff = 1'h0;
  end
  if (reset) begin
    ifc_dma_access_ok_prev = 1'h0;
  end
  if (reset) begin
    iccm_ecc_corr_data_ff = 39'h0;
  end
  if (reset) begin
    dma_mem_addr_ff = 2'h0;
  end
  if (reset) begin
    dma_mem_tag_ff = 3'h0;
  end
  if (reset) begin
    iccm_dma_rtag_temp = 3'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_temp = 1'h0;
  end
  if (reset) begin
    iccm_dma_ecc_error = 1'h0;
  end
  if (reset) begin
    iccm_dma_rdata_temp = 64'h0;
  end
  if (reset) begin
    iccm_ecc_corr_index_ff = 14'h0;
  end
  if (reset) begin
    iccm_rd_ecc_single_err_ff = 1'h0;
  end
  if (reset) begin
    iccm_rw_addr_f = 14'h0;
  end
  if (reset) begin
    ifu_status_wr_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_wr_en_ff = 1'h0;
  end
  if (reset) begin
    way_status_new_ff = 1'h0;
  end
  if (reset) begin
    ifu_tag_wren_ff = 2'h0;
  end
  if (reset) begin
    ic_valid_ff = 1'h0;
  end
  if (reset) begin
    _T_9748 = 1'h0;
  end
  if (reset) begin
    _T_9749 = 1'h0;
  end
  if (reset) begin
    _T_9750 = 1'h0;
  end
  if (reset) begin
    _T_9754 = 1'h0;
  end
  if (reset) begin
    _T_9755 = 1'h0;
  end
  if (reset) begin
    _T_9776 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_2_io_l1clk) begin
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge io_free_clk) begin
    reset_ic_ff <= _T_298 & _T_299;
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= _T_317 & _T_318;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= _T_22 & _T_319;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2660 & _T_2664;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2451) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2453) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2463) begin
        perr_state <= 3'h0;
      end else if (_T_2466) begin
        if (_T_2469) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2473) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2477) begin
        err_stop_state <= 2'h1;
      end else if (_T_2482) begin
        if (_T_2484) begin
          err_stop_state <= 2'h0;
        end else if (_T_2505) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2509) begin
        if (_T_2484) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2526) begin
        if (_T_2530) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf | ifc_region_acc_fault_memory_bf;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= _T_2582 | _T_2583;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= {_T_1353,ic_miss_buff_data_valid_in_0};
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= _T_2590 | _T_2592;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= _T_334 | reset_tag_valid_for_miss;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_3946) begin
      ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_ic_rw_int_addr_ff <= ifu_ic_rw_int_addr[11:5];
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_0 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_1 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_2 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_3 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_4 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_5 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_6 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_7 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_8 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_9 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_10 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_11 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_12 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_13 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_14 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_15 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_16 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_17 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_18 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_19 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_20 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_21 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_22 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_23 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_24 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_25 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_26 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_27 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_28 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_29 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_30 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_31 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_32 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_33 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_34 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_35 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_36 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_37 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_38 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_39 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_40 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_41 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_42 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_43 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_44 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_45 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_46 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_47 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_48 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_49 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_50 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_51 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_52 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_53 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_54 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_55 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_56 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_57 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_58 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_59 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_60 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_61 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_62 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_63 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_64 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_65 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_66 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_67 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_68 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_69 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_70 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_71 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_72 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_73 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_74 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_75 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_76 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_77 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_78 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_79 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_80 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_81 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_82 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_83 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_84 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_85 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_86 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_87 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_88 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_89 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_90 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_91 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_92 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_93 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_94 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_95 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_96 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_97 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_98 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_99 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_100 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_101 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_102 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_103 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_104 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_105 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_106 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_107 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_108 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_109 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_110 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_111 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_112 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_113 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_114 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_115 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_116 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_117 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_118 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_119 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_3970) begin
      way_status_out_120 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_3974) begin
      way_status_out_121 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_3978) begin
      way_status_out_122 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_123 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_124 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_3990) begin
      way_status_out_125 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_3994) begin
      way_status_out_126 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_3998) begin
      way_status_out_127 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      tagv_mb_scnd_ff <= 2'h0;
    end else if (!(_T_19)) begin
      tagv_mb_scnd_ff <= _T_198;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err_data & _T_2578;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_290;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= _T_295;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_231) begin
      bus_rd_addr_count <= imb_ff[4:2];
    end else if (scnd_miss_req_q) begin
      bus_rd_addr_count <= imb_scnd_ff[4:2];
    end else if (bus_cmd_sent) begin
      bus_rd_addr_count <= _T_2598;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= _T_233 & _T_209;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= _T_1509 | _T_1514;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= {_T_1393,ic_miss_buff_data_error_in_0};
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else begin
      ic_debug_ict_array_sel_ff <= io_ic_debug_rd_en & io_ic_debug_tag_array;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5591) begin
      ic_tag_valid_out_1_0 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5606) begin
      ic_tag_valid_out_1_1 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5621) begin
      ic_tag_valid_out_1_2 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5636) begin
      ic_tag_valid_out_1_3 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5651) begin
      ic_tag_valid_out_1_4 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5666) begin
      ic_tag_valid_out_1_5 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5681) begin
      ic_tag_valid_out_1_6 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5696) begin
      ic_tag_valid_out_1_7 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5711) begin
      ic_tag_valid_out_1_8 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5726) begin
      ic_tag_valid_out_1_9 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5741) begin
      ic_tag_valid_out_1_10 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5756) begin
      ic_tag_valid_out_1_11 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5771) begin
      ic_tag_valid_out_1_12 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5786) begin
      ic_tag_valid_out_1_13 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5801) begin
      ic_tag_valid_out_1_14 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5816) begin
      ic_tag_valid_out_1_15 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5831) begin
      ic_tag_valid_out_1_16 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5846) begin
      ic_tag_valid_out_1_17 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5861) begin
      ic_tag_valid_out_1_18 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5876) begin
      ic_tag_valid_out_1_19 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5891) begin
      ic_tag_valid_out_1_20 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5906) begin
      ic_tag_valid_out_1_21 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5921) begin
      ic_tag_valid_out_1_22 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5936) begin
      ic_tag_valid_out_1_23 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_5951) begin
      ic_tag_valid_out_1_24 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_5966) begin
      ic_tag_valid_out_1_25 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_5981) begin
      ic_tag_valid_out_1_26 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_5996) begin
      ic_tag_valid_out_1_27 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6011) begin
      ic_tag_valid_out_1_28 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6026) begin
      ic_tag_valid_out_1_29 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6041) begin
      ic_tag_valid_out_1_30 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6056) begin
      ic_tag_valid_out_1_31 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6551) begin
      ic_tag_valid_out_1_32 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6566) begin
      ic_tag_valid_out_1_33 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6581) begin
      ic_tag_valid_out_1_34 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6596) begin
      ic_tag_valid_out_1_35 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6611) begin
      ic_tag_valid_out_1_36 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6626) begin
      ic_tag_valid_out_1_37 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6641) begin
      ic_tag_valid_out_1_38 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6656) begin
      ic_tag_valid_out_1_39 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6671) begin
      ic_tag_valid_out_1_40 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6686) begin
      ic_tag_valid_out_1_41 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6701) begin
      ic_tag_valid_out_1_42 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6716) begin
      ic_tag_valid_out_1_43 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6731) begin
      ic_tag_valid_out_1_44 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6746) begin
      ic_tag_valid_out_1_45 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6761) begin
      ic_tag_valid_out_1_46 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6776) begin
      ic_tag_valid_out_1_47 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6791) begin
      ic_tag_valid_out_1_48 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6806) begin
      ic_tag_valid_out_1_49 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6821) begin
      ic_tag_valid_out_1_50 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6836) begin
      ic_tag_valid_out_1_51 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6851) begin
      ic_tag_valid_out_1_52 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6866) begin
      ic_tag_valid_out_1_53 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6881) begin
      ic_tag_valid_out_1_54 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6896) begin
      ic_tag_valid_out_1_55 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6911) begin
      ic_tag_valid_out_1_56 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6926) begin
      ic_tag_valid_out_1_57 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6941) begin
      ic_tag_valid_out_1_58 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_6956) begin
      ic_tag_valid_out_1_59 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_6971) begin
      ic_tag_valid_out_1_60 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_6986) begin
      ic_tag_valid_out_1_61 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7001) begin
      ic_tag_valid_out_1_62 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7016) begin
      ic_tag_valid_out_1_63 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7511) begin
      ic_tag_valid_out_1_64 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7526) begin
      ic_tag_valid_out_1_65 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7541) begin
      ic_tag_valid_out_1_66 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7556) begin
      ic_tag_valid_out_1_67 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7571) begin
      ic_tag_valid_out_1_68 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7586) begin
      ic_tag_valid_out_1_69 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7601) begin
      ic_tag_valid_out_1_70 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7616) begin
      ic_tag_valid_out_1_71 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7631) begin
      ic_tag_valid_out_1_72 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7646) begin
      ic_tag_valid_out_1_73 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7661) begin
      ic_tag_valid_out_1_74 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7676) begin
      ic_tag_valid_out_1_75 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7691) begin
      ic_tag_valid_out_1_76 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7706) begin
      ic_tag_valid_out_1_77 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7721) begin
      ic_tag_valid_out_1_78 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7736) begin
      ic_tag_valid_out_1_79 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7751) begin
      ic_tag_valid_out_1_80 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7766) begin
      ic_tag_valid_out_1_81 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7781) begin
      ic_tag_valid_out_1_82 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7796) begin
      ic_tag_valid_out_1_83 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7811) begin
      ic_tag_valid_out_1_84 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7826) begin
      ic_tag_valid_out_1_85 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7841) begin
      ic_tag_valid_out_1_86 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7856) begin
      ic_tag_valid_out_1_87 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7871) begin
      ic_tag_valid_out_1_88 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7886) begin
      ic_tag_valid_out_1_89 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7901) begin
      ic_tag_valid_out_1_90 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7916) begin
      ic_tag_valid_out_1_91 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7931) begin
      ic_tag_valid_out_1_92 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7946) begin
      ic_tag_valid_out_1_93 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_7961) begin
      ic_tag_valid_out_1_94 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_7976) begin
      ic_tag_valid_out_1_95 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8471) begin
      ic_tag_valid_out_1_96 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8486) begin
      ic_tag_valid_out_1_97 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8501) begin
      ic_tag_valid_out_1_98 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8516) begin
      ic_tag_valid_out_1_99 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8531) begin
      ic_tag_valid_out_1_100 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8546) begin
      ic_tag_valid_out_1_101 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8561) begin
      ic_tag_valid_out_1_102 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8576) begin
      ic_tag_valid_out_1_103 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8591) begin
      ic_tag_valid_out_1_104 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8606) begin
      ic_tag_valid_out_1_105 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8621) begin
      ic_tag_valid_out_1_106 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8636) begin
      ic_tag_valid_out_1_107 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8651) begin
      ic_tag_valid_out_1_108 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8666) begin
      ic_tag_valid_out_1_109 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8681) begin
      ic_tag_valid_out_1_110 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8696) begin
      ic_tag_valid_out_1_111 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8711) begin
      ic_tag_valid_out_1_112 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8726) begin
      ic_tag_valid_out_1_113 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8741) begin
      ic_tag_valid_out_1_114 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8756) begin
      ic_tag_valid_out_1_115 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8771) begin
      ic_tag_valid_out_1_116 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8786) begin
      ic_tag_valid_out_1_117 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8801) begin
      ic_tag_valid_out_1_118 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8816) begin
      ic_tag_valid_out_1_119 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8831) begin
      ic_tag_valid_out_1_120 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8846) begin
      ic_tag_valid_out_1_121 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8861) begin
      ic_tag_valid_out_1_122 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8876) begin
      ic_tag_valid_out_1_123 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8891) begin
      ic_tag_valid_out_1_124 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8906) begin
      ic_tag_valid_out_1_125 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8921) begin
      ic_tag_valid_out_1_126 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8936) begin
      ic_tag_valid_out_1_127 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5111) begin
      ic_tag_valid_out_0_0 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5126) begin
      ic_tag_valid_out_0_1 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5141) begin
      ic_tag_valid_out_0_2 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5156) begin
      ic_tag_valid_out_0_3 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5171) begin
      ic_tag_valid_out_0_4 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5186) begin
      ic_tag_valid_out_0_5 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5201) begin
      ic_tag_valid_out_0_6 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5216) begin
      ic_tag_valid_out_0_7 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5231) begin
      ic_tag_valid_out_0_8 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5246) begin
      ic_tag_valid_out_0_9 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5261) begin
      ic_tag_valid_out_0_10 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5276) begin
      ic_tag_valid_out_0_11 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5291) begin
      ic_tag_valid_out_0_12 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5306) begin
      ic_tag_valid_out_0_13 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5321) begin
      ic_tag_valid_out_0_14 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5336) begin
      ic_tag_valid_out_0_15 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5351) begin
      ic_tag_valid_out_0_16 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5366) begin
      ic_tag_valid_out_0_17 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5381) begin
      ic_tag_valid_out_0_18 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5396) begin
      ic_tag_valid_out_0_19 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5411) begin
      ic_tag_valid_out_0_20 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5426) begin
      ic_tag_valid_out_0_21 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5441) begin
      ic_tag_valid_out_0_22 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5456) begin
      ic_tag_valid_out_0_23 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5471) begin
      ic_tag_valid_out_0_24 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5486) begin
      ic_tag_valid_out_0_25 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5501) begin
      ic_tag_valid_out_0_26 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5516) begin
      ic_tag_valid_out_0_27 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5531) begin
      ic_tag_valid_out_0_28 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5546) begin
      ic_tag_valid_out_0_29 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5561) begin
      ic_tag_valid_out_0_30 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5576) begin
      ic_tag_valid_out_0_31 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6071) begin
      ic_tag_valid_out_0_32 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6086) begin
      ic_tag_valid_out_0_33 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6101) begin
      ic_tag_valid_out_0_34 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6116) begin
      ic_tag_valid_out_0_35 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6131) begin
      ic_tag_valid_out_0_36 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6146) begin
      ic_tag_valid_out_0_37 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6161) begin
      ic_tag_valid_out_0_38 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6176) begin
      ic_tag_valid_out_0_39 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6191) begin
      ic_tag_valid_out_0_40 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6206) begin
      ic_tag_valid_out_0_41 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6221) begin
      ic_tag_valid_out_0_42 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6236) begin
      ic_tag_valid_out_0_43 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6251) begin
      ic_tag_valid_out_0_44 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6266) begin
      ic_tag_valid_out_0_45 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6281) begin
      ic_tag_valid_out_0_46 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6296) begin
      ic_tag_valid_out_0_47 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6311) begin
      ic_tag_valid_out_0_48 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6326) begin
      ic_tag_valid_out_0_49 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6341) begin
      ic_tag_valid_out_0_50 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6356) begin
      ic_tag_valid_out_0_51 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6371) begin
      ic_tag_valid_out_0_52 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6386) begin
      ic_tag_valid_out_0_53 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6401) begin
      ic_tag_valid_out_0_54 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6416) begin
      ic_tag_valid_out_0_55 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6431) begin
      ic_tag_valid_out_0_56 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6446) begin
      ic_tag_valid_out_0_57 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6461) begin
      ic_tag_valid_out_0_58 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6476) begin
      ic_tag_valid_out_0_59 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6491) begin
      ic_tag_valid_out_0_60 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6506) begin
      ic_tag_valid_out_0_61 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6521) begin
      ic_tag_valid_out_0_62 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6536) begin
      ic_tag_valid_out_0_63 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7031) begin
      ic_tag_valid_out_0_64 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7046) begin
      ic_tag_valid_out_0_65 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7061) begin
      ic_tag_valid_out_0_66 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7076) begin
      ic_tag_valid_out_0_67 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7091) begin
      ic_tag_valid_out_0_68 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7106) begin
      ic_tag_valid_out_0_69 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7121) begin
      ic_tag_valid_out_0_70 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7136) begin
      ic_tag_valid_out_0_71 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7151) begin
      ic_tag_valid_out_0_72 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7166) begin
      ic_tag_valid_out_0_73 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7181) begin
      ic_tag_valid_out_0_74 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7196) begin
      ic_tag_valid_out_0_75 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7211) begin
      ic_tag_valid_out_0_76 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7226) begin
      ic_tag_valid_out_0_77 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7241) begin
      ic_tag_valid_out_0_78 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7256) begin
      ic_tag_valid_out_0_79 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7271) begin
      ic_tag_valid_out_0_80 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7286) begin
      ic_tag_valid_out_0_81 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7301) begin
      ic_tag_valid_out_0_82 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7316) begin
      ic_tag_valid_out_0_83 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7331) begin
      ic_tag_valid_out_0_84 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7346) begin
      ic_tag_valid_out_0_85 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7361) begin
      ic_tag_valid_out_0_86 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7376) begin
      ic_tag_valid_out_0_87 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7391) begin
      ic_tag_valid_out_0_88 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7406) begin
      ic_tag_valid_out_0_89 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7421) begin
      ic_tag_valid_out_0_90 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7436) begin
      ic_tag_valid_out_0_91 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7451) begin
      ic_tag_valid_out_0_92 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7466) begin
      ic_tag_valid_out_0_93 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7481) begin
      ic_tag_valid_out_0_94 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7496) begin
      ic_tag_valid_out_0_95 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_7991) begin
      ic_tag_valid_out_0_96 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8006) begin
      ic_tag_valid_out_0_97 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8021) begin
      ic_tag_valid_out_0_98 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8036) begin
      ic_tag_valid_out_0_99 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8051) begin
      ic_tag_valid_out_0_100 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8066) begin
      ic_tag_valid_out_0_101 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8081) begin
      ic_tag_valid_out_0_102 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8096) begin
      ic_tag_valid_out_0_103 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8111) begin
      ic_tag_valid_out_0_104 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8126) begin
      ic_tag_valid_out_0_105 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8141) begin
      ic_tag_valid_out_0_106 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8156) begin
      ic_tag_valid_out_0_107 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8171) begin
      ic_tag_valid_out_0_108 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8186) begin
      ic_tag_valid_out_0_109 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8201) begin
      ic_tag_valid_out_0_110 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8216) begin
      ic_tag_valid_out_0_111 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8231) begin
      ic_tag_valid_out_0_112 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8246) begin
      ic_tag_valid_out_0_113 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8261) begin
      ic_tag_valid_out_0_114 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8276) begin
      ic_tag_valid_out_0_115 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8291) begin
      ic_tag_valid_out_0_116 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8306) begin
      ic_tag_valid_out_0_117 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8321) begin
      ic_tag_valid_out_0_118 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8336) begin
      ic_tag_valid_out_0_119 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8351) begin
      ic_tag_valid_out_0_120 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8366) begin
      ic_tag_valid_out_0_121 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8381) begin
      ic_tag_valid_out_0_122 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8396) begin
      ic_tag_valid_out_0_123 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8411) begin
      ic_tag_valid_out_0_124 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8426) begin
      ic_tag_valid_out_0_125 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8441) begin
      ic_tag_valid_out_0_126 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8456) begin
      ic_tag_valid_out_0_127 <= _T_5103;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_1211 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1211 <= _T_1210;
    end else begin
      _T_1211 <= io_ic_debug_rd_data;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_memory_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_memory_f <= _T_9835 & io_ifc_fetch_req_bf;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= perr_state == 3'h4;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_cmd_req_hold <= 1'h0;
    end else begin
      bus_cmd_req_hold <= _T_2555 & _T_2574;
    end
  end
  always @(posedge rvclkhdr_69_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else begin
      ifu_bus_cmd_valid <= _T_2545 & _T_2551;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (bus_cmd_beat_en) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= _T_2650 & _T_2651;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3881;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rtag_temp <= 3'h0;
    end else begin
      iccm_dma_rtag_temp <= dma_mem_tag_ff;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_temp <= 1'h0;
    end else begin
      iccm_dma_rvalid_temp <= iccm_dma_rvalid_in;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_ecc_error <= 1'h0;
    end else begin
      iccm_dma_ecc_error <= |iccm_double_ecc_error;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rdata_temp <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata_temp <= _T_3055;
    end else begin
      iccm_dma_rdata_temp <= _T_3056;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3877;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= _T_3872 & _T_319;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3946) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en | _T_3949;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_3949) begin
      way_status_new_ff <= io_ic_debug_wr_data[4];
    end else if (_T_9726) begin
      way_status_new_ff <= replace_way_mb_any_0;
    end else begin
      way_status_new_ff <= way_status_hit_new;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren | ic_debug_tag_wr_en;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3949) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9748 <= 1'h0;
    end else begin
      _T_9748 <= _T_233 & _T_209;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9749 <= 1'h0;
    end else begin
      _T_9749 <= _T_225 & _T_247;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9750 <= 1'h0;
    end else begin
      _T_9750 <= ic_byp_hit_f & ifu_byp_data_err_new;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9754 <= 1'h0;
    end else begin
      _T_9754 <= _T_9752 & miss_pending;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9755 <= 1'h0;
    end else begin
      _T_9755 <= _T_2569 & _T_2574;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_9776 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_9776 <= ic_debug_rd_en_ff;
    end
  end
endmodule
