module el2_ifu_compress_ctl(
  input         clock,
  input         reset,
  input  [15:0] io_in,
  output [31:0] io_out
);
  wire  _T_1 = io_in[1:0] != 2'h3; // @[el2_ifu_compress_ctl.scala 192:26]
  wire [31:0] _T_3 = {16'h0,io_in}; // @[Cat.scala 29:58]
  wire  _T_5 = |_T_3[12:5]; // @[el2_ifu_compress_ctl.scala 48:29]
  wire [6:0] _T_6 = _T_5 ? 7'h13 : 7'h1f; // @[el2_ifu_compress_ctl.scala 48:20]
  wire [29:0] _T_20 = {_T_3[10:7],_T_3[12:11],_T_3[5],_T_3[6],2'h0,5'h2,3'h0,2'h1,_T_3[4:2],_T_6}; // @[Cat.scala 29:58]
  wire [7:0] _T_30 = {_T_3[6:5],_T_3[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [27:0] _T_38 = {_T_3[6:5],_T_3[12:10],3'h0,2'h1,_T_3[9:7],3'h3,2'h1,_T_3[4:2],7'h7}; // @[Cat.scala 29:58]
  wire [6:0] _T_52 = {_T_3[5],_T_3[12:10],_T_3[6],2'h0}; // @[Cat.scala 29:58]
  wire [26:0] _T_60 = {_T_3[5],_T_3[12:10],_T_3[6],2'h0,2'h1,_T_3[9:7],3'h2,2'h1,_T_3[4:2],7'h3}; // @[Cat.scala 29:58]
  wire [27:0] _T_80 = {_T_3[6:5],_T_3[12:10],3'h0,2'h1,_T_3[9:7],3'h3,2'h1,_T_3[4:2],7'h3}; // @[Cat.scala 29:58]
  wire [26:0] _T_111 = {_T_52[6:5],2'h1,_T_3[4:2],2'h1,_T_3[9:7],3'h2,_T_52[4:0],7'h3f}; // @[Cat.scala 29:58]
  wire [27:0] _T_138 = {_T_30[7:5],2'h1,_T_3[4:2],2'h1,_T_3[9:7],3'h3,_T_30[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [26:0] _T_169 = {_T_52[6:5],2'h1,_T_3[4:2],2'h1,_T_3[9:7],3'h2,_T_52[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [27:0] _T_196 = {_T_30[7:5],2'h1,_T_3[4:2],2'h1,_T_3[9:7],3'h3,_T_30[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [6:0] _T_207 = _T_3[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_209 = {_T_207,_T_3[6:2]}; // @[Cat.scala 29:58]
  wire [31:0] _T_215 = {_T_207,_T_3[6:2],_T_3[11:7],3'h0,_T_3[11:7],7'h13}; // @[Cat.scala 29:58]
  wire  _T_223 = |_T_3[11:7]; // @[el2_ifu_compress_ctl.scala 72:24]
  wire [6:0] _T_224 = _T_223 ? 7'h1b : 7'h1f; // @[el2_ifu_compress_ctl.scala 72:20]
  wire [31:0] _T_235 = {_T_207,_T_3[6:2],_T_3[11:7],3'h0,_T_3[11:7],_T_224}; // @[Cat.scala 29:58]
  wire [31:0] _T_251 = {_T_207,_T_3[6:2],5'h0,3'h0,_T_3[11:7],7'h13}; // @[Cat.scala 29:58]
  wire  _T_262 = |_T_209; // @[el2_ifu_compress_ctl.scala 85:29]
  wire [6:0] _T_263 = _T_262 ? 7'h37 : 7'h3f; // @[el2_ifu_compress_ctl.scala 85:20]
  wire [14:0] _T_266 = _T_3[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_269 = {_T_266,_T_3[6:2],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_273 = {_T_269[31:12],_T_3[11:7],_T_263}; // @[Cat.scala 29:58]
  wire  _T_281 = _T_3[11:7] == 5'h0; // @[el2_ifu_compress_ctl.scala 87:14]
  wire  _T_283 = _T_3[11:7] == 5'h2; // @[el2_ifu_compress_ctl.scala 87:27]
  wire  _T_284 = _T_281 | _T_283; // @[el2_ifu_compress_ctl.scala 87:21]
  wire [6:0] _T_291 = _T_262 ? 7'h13 : 7'h1f; // @[el2_ifu_compress_ctl.scala 81:20]
  wire [2:0] _T_294 = _T_3[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_309 = {_T_294,_T_3[4:3],_T_3[5],_T_3[2],_T_3[6],4'h0,_T_3[11:7],3'h0,_T_3[11:7],_T_291}; // @[Cat.scala 29:58]
  wire [31:0] _T_316_bits = _T_284 ? _T_309 : _T_273; // @[el2_ifu_compress_ctl.scala 87:10]
  wire [25:0] _T_327 = {_T_3[12],_T_3[6:2],2'h1,_T_3[9:7],3'h5,2'h1,_T_3[9:7],7'h13}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_172 = {{5'd0}, _T_327}; // @[el2_ifu_compress_ctl.scala 94:23]
  wire [30:0] _T_339 = _GEN_172 | 31'h40000000; // @[el2_ifu_compress_ctl.scala 94:23]
  wire [31:0] _T_352 = {_T_207,_T_3[6:2],2'h1,_T_3[9:7],3'h7,2'h1,_T_3[9:7],7'h13}; // @[Cat.scala 29:58]
  wire [2:0] _T_356 = {_T_3[12],_T_3[6:5]}; // @[Cat.scala 29:58]
  wire  _T_358 = _T_3[6:5] == 2'h0; // @[el2_ifu_compress_ctl.scala 98:30]
  wire [30:0] _T_359 = _T_358 ? 31'h40000000 : 31'h0; // @[el2_ifu_compress_ctl.scala 98:22]
  wire [6:0] _T_361 = _T_3[12] ? 7'h3b : 7'h33; // @[el2_ifu_compress_ctl.scala 99:22]
  wire [2:0] _GEN_1 = 3'h1 == _T_356 ? 3'h4 : 3'h0; // @[Cat.scala 29:58]
  wire [2:0] _GEN_2 = 3'h2 == _T_356 ? 3'h6 : _GEN_1; // @[Cat.scala 29:58]
  wire [2:0] _GEN_3 = 3'h3 == _T_356 ? 3'h7 : _GEN_2; // @[Cat.scala 29:58]
  wire [2:0] _GEN_4 = 3'h4 == _T_356 ? 3'h0 : _GEN_3; // @[Cat.scala 29:58]
  wire [2:0] _GEN_5 = 3'h5 == _T_356 ? 3'h0 : _GEN_4; // @[Cat.scala 29:58]
  wire [2:0] _GEN_6 = 3'h6 == _T_356 ? 3'h2 : _GEN_5; // @[Cat.scala 29:58]
  wire [2:0] _GEN_7 = 3'h7 == _T_356 ? 3'h3 : _GEN_6; // @[Cat.scala 29:58]
  wire [24:0] _T_371 = {2'h1,_T_3[4:2],2'h1,_T_3[9:7],_GEN_7,2'h1,_T_3[9:7],_T_361}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_173 = {{6'd0}, _T_371}; // @[el2_ifu_compress_ctl.scala 100:43]
  wire [30:0] _T_372 = _GEN_173 | _T_359; // @[el2_ifu_compress_ctl.scala 100:43]
  wire [31:0] _T_373_0 = {{6'd0}, _T_327}; // @[el2_ifu_compress_ctl.scala 102:19 el2_ifu_compress_ctl.scala 102:19]
  wire [31:0] _T_373_1 = {{1'd0}, _T_339}; // @[el2_ifu_compress_ctl.scala 102:19 el2_ifu_compress_ctl.scala 102:19]
  wire [31:0] _GEN_9 = 2'h1 == _T_3[11:10] ? _T_373_1 : _T_373_0; // @[el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_10 = 2'h2 == _T_3[11:10] ? _T_352 : _GEN_9; // @[el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _T_373_3 = {{1'd0}, _T_372}; // @[el2_ifu_compress_ctl.scala 102:19 el2_ifu_compress_ctl.scala 102:19]
  wire [31:0] _GEN_11 = 2'h3 == _T_3[11:10] ? _T_373_3 : _GEN_10; // @[el2_ifu_compress_ctl.scala 17:14]
  wire [9:0] _T_385 = _T_3[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  wire [20:0] _T_400 = {_T_385,_T_3[8],_T_3[10:9],_T_3[6],_T_3[7],_T_3[2],_T_3[11],_T_3[5:3],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_463 = {_T_400[20],_T_400[10:1],_T_400[11],_T_400[19:12],5'h0,7'h6f}; // @[Cat.scala 29:58]
  wire [4:0] _T_472 = _T_3[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [12:0] _T_481 = {_T_472,_T_3[6:5],_T_3[2],_T_3[11:10],_T_3[4:3],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_530 = {_T_481[12],_T_481[10:5],5'h0,2'h1,_T_3[9:7],3'h0,_T_481[4:1],_T_481[11],7'h63}; // @[Cat.scala 29:58]
  wire [31:0] _T_597 = {_T_481[12],_T_481[10:5],5'h0,2'h1,_T_3[9:7],3'h1,_T_481[4:1],_T_481[11],7'h63}; // @[Cat.scala 29:58]
  wire [6:0] _T_604 = _T_223 ? 7'h3 : 7'h1f; // @[el2_ifu_compress_ctl.scala 108:23]
  wire [25:0] _T_613 = {_T_3[12],_T_3[6:2],_T_3[11:7],3'h1,_T_3[11:7],7'h13}; // @[Cat.scala 29:58]
  wire [28:0] _T_629 = {_T_3[4:2],_T_3[12],_T_3[6:5],3'h0,5'h2,3'h3,_T_3[11:7],7'h7}; // @[Cat.scala 29:58]
  wire [27:0] _T_644 = {_T_3[3:2],_T_3[12],_T_3[6:4],2'h0,5'h2,3'h2,_T_3[11:7],_T_604}; // @[Cat.scala 29:58]
  wire [28:0] _T_659 = {_T_3[4:2],_T_3[12],_T_3[6:5],3'h0,5'h2,3'h3,_T_3[11:7],_T_604}; // @[Cat.scala 29:58]
  wire [24:0] _T_669 = {_T_3[6:2],5'h0,3'h0,_T_3[11:7],7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _T_680 = {_T_3[6:2],_T_3[11:7],3'h0,_T_3[11:7],7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _T_691 = {_T_3[6:2],_T_3[11:7],3'h0,12'h67}; // @[Cat.scala 29:58]
  wire [24:0] _T_693 = {_T_691[24:7],7'h1f}; // @[Cat.scala 29:58]
  wire [24:0] _T_696 = _T_223 ? _T_691 : _T_693; // @[el2_ifu_compress_ctl.scala 129:33]
  wire  _T_702 = |_T_3[6:2]; // @[el2_ifu_compress_ctl.scala 130:27]
  wire [31:0] _T_673_bits = {{7'd0}, _T_669}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _T_700_bits = {{7'd0}, _T_696}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _T_703_bits = _T_702 ? _T_673_bits : _T_700_bits; // @[el2_ifu_compress_ctl.scala 130:22]
  wire [24:0] _T_709 = {_T_3[6:2],_T_3[11:7],3'h0,12'he7}; // @[Cat.scala 29:58]
  wire [24:0] _T_711 = {_T_691[24:7],7'h73}; // @[Cat.scala 29:58]
  wire [24:0] _T_712 = _T_711 | 25'h100000; // @[el2_ifu_compress_ctl.scala 132:46]
  wire [24:0] _T_715 = _T_223 ? _T_709 : _T_712; // @[el2_ifu_compress_ctl.scala 133:33]
  wire [31:0] _T_685_bits = {{7'd0}, _T_680}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _T_719_bits = {{7'd0}, _T_715}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _T_722_bits = _T_702 ? _T_685_bits : _T_719_bits; // @[el2_ifu_compress_ctl.scala 134:25]
  wire [31:0] _T_724_bits = _T_3[12] ? _T_722_bits : _T_703_bits; // @[el2_ifu_compress_ctl.scala 135:10]
  wire [8:0] _T_728 = {_T_3[9:7],_T_3[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [28:0] _T_740 = {_T_728[8:5],_T_3[6:2],5'h2,3'h3,_T_728[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [7:0] _T_748 = {_T_3[8:7],_T_3[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [27:0] _T_760 = {_T_748[7:5],_T_3[6:2],5'h2,3'h2,_T_748[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [28:0] _T_780 = {_T_728[8:5],_T_3[6:2],5'h2,3'h3,_T_728[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [4:0] _T_828 = {_T_3[1:0],_T_3[15:13]}; // @[Cat.scala 29:58]
  wire [31:0] _T_26_bits = {{2'd0}, _T_20}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _T_46_bits = {{4'd0}, _T_38}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_17 = 5'h1 == _T_828 ? _T_46_bits : _T_26_bits; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_68_bits = {{5'd0}, _T_60}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_22 = 5'h2 == _T_828 ? _T_68_bits : _GEN_17; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_88_bits = {{4'd0}, _T_80}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_27 = 5'h3 == _T_828 ? _T_88_bits : _GEN_22; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_119_bits = {{5'd0}, _T_111}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_32 = 5'h4 == _T_828 ? _T_119_bits : _GEN_27; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_146_bits = {{4'd0}, _T_138}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_37 = 5'h5 == _T_828 ? _T_146_bits : _GEN_32; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_177_bits = {{5'd0}, _T_169}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_42 = 5'h6 == _T_828 ? _T_177_bits : _GEN_37; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_204_bits = {{4'd0}, _T_196}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_47 = 5'h7 == _T_828 ? _T_204_bits : _GEN_42; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_52 = 5'h8 == _T_828 ? _T_215 : _GEN_47; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_57 = 5'h9 == _T_828 ? _T_235 : _GEN_52; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_62 = 5'ha == _T_828 ? _T_251 : _GEN_57; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_67 = 5'hb == _T_828 ? _T_316_bits : _GEN_62; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_72 = 5'hc == _T_828 ? _GEN_11 : _GEN_67; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_77 = 5'hd == _T_828 ? _T_463 : _GEN_72; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_82 = 5'he == _T_828 ? _T_530 : _GEN_77; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_87 = 5'hf == _T_828 ? _T_597 : _GEN_82; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_618_bits = {{6'd0}, _T_613}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_92 = 5'h10 == _T_828 ? _T_618_bits : _GEN_87; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_633_bits = {{3'd0}, _T_629}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_97 = 5'h11 == _T_828 ? _T_633_bits : _GEN_92; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_648_bits = {{4'd0}, _T_644}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_102 = 5'h12 == _T_828 ? _T_648_bits : _GEN_97; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_663_bits = {{3'd0}, _T_659}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_107 = 5'h13 == _T_828 ? _T_663_bits : _GEN_102; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_112 = 5'h14 == _T_828 ? _T_724_bits : _GEN_107; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_744_bits = {{3'd0}, _T_740}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_117 = 5'h15 == _T_828 ? _T_744_bits : _GEN_112; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_764_bits = {{4'd0}, _T_760}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_122 = 5'h16 == _T_828 ? _T_764_bits : _GEN_117; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _T_784_bits = {{3'd0}, _T_780}; // @[el2_ifu_compress_ctl.scala 16:19 el2_ifu_compress_ctl.scala 17:14]
  wire [31:0] _GEN_127 = 5'h17 == _T_828 ? _T_784_bits : _GEN_122; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_132 = 5'h18 == _T_828 ? _T_3 : _GEN_127; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_137 = 5'h19 == _T_828 ? _T_3 : _GEN_132; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_142 = 5'h1a == _T_828 ? _T_3 : _GEN_137; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_147 = 5'h1b == _T_828 ? _T_3 : _GEN_142; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_152 = 5'h1c == _T_828 ? _T_3 : _GEN_147; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_157 = 5'h1d == _T_828 ? _T_3 : _GEN_152; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_162 = 5'h1e == _T_828 ? _T_3 : _GEN_157; // @[el2_ifu_compress_ctl.scala 195:18]
  wire [31:0] _GEN_167 = 5'h1f == _T_828 ? _T_3 : _GEN_162; // @[el2_ifu_compress_ctl.scala 195:18]
  assign io_out = _T_1 ? 32'h0 : _GEN_167; // @[el2_ifu_compress_ctl.scala 195:12]
endmodule
