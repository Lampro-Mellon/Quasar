module rvclkhdr(
  input   io_clk,
  input   io_en
);
  wire  clkhdr_Q; // @[lib.scala 334:26]
  wire  clkhdr_CK; // @[lib.scala 334:26]
  wire  clkhdr_EN; // @[lib.scala 334:26]
  wire  clkhdr_SE; // @[lib.scala 334:26]
  gated_latch clkhdr ( // @[lib.scala 334:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign clkhdr_CK = io_clk; // @[lib.scala 336:18]
  assign clkhdr_EN = io_en; // @[lib.scala 337:18]
  assign clkhdr_SE = 1'h0; // @[lib.scala 338:18]
endmodule
module ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_l2clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_mem_ctrl_dec_tlu_flush_err_wb,
  input         io_dec_mem_ctrl_dec_tlu_i0_commit_cmt,
  input         io_dec_mem_ctrl_dec_tlu_force_halt,
  input         io_dec_mem_ctrl_dec_tlu_fence_i_wb,
  input  [70:0] io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid,
  input         io_dec_mem_ctrl_dec_tlu_core_ecc_disable,
  output        io_dec_mem_ctrl_ifu_pmu_ic_miss,
  output        io_dec_mem_ctrl_ifu_pmu_ic_hit,
  output        io_dec_mem_ctrl_ifu_pmu_bus_error,
  output        io_dec_mem_ctrl_ifu_pmu_bus_busy,
  output        io_dec_mem_ctrl_ifu_pmu_bus_trxn,
  output        io_dec_mem_ctrl_ifu_ic_error_start,
  output        io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err,
  output [70:0] io_dec_mem_ctrl_ifu_ic_debug_rd_data,
  output        io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid,
  output        io_dec_mem_ctrl_ifu_miss_state_idle,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_ar_ready,
  output        io_ifu_axi_ar_valid,
  output [2:0]  io_ifu_axi_ar_bits_id,
  output [31:0] io_ifu_axi_ar_bits_addr,
  output [3:0]  io_ifu_axi_ar_bits_region,
  output        io_ifu_axi_r_ready,
  input         io_ifu_axi_r_valid,
  input  [2:0]  io_ifu_axi_r_bits_id,
  input  [63:0] io_ifu_axi_r_bits_data,
  input  [1:0]  io_ifu_axi_r_bits_resp,
  input         io_ifu_bus_clk_en,
  input         io_dma_mem_ctl_dma_iccm_req,
  input  [31:0] io_dma_mem_ctl_dma_mem_addr,
  input  [2:0]  io_dma_mem_ctl_dma_mem_sz,
  input         io_dma_mem_ctl_dma_mem_write,
  input  [63:0] io_dma_mem_ctl_dma_mem_wdata,
  input  [2:0]  io_dma_mem_ctl_dma_mem_tag,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [2:0]  io_iccm_wr_size,
  output [77:0] io_iccm_wr_data,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_tag_valid,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [9:0]  io_ic_debug_addr,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ic_tag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input  [1:0]  io_ifu_fetch_val,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  input         io_dec_tlu_flush_lower_wb,
  output [1:0]  io_iccm_rd_ecc_double_err,
  output        io_iccm_dma_sb_error,
  output        io_ic_hit_f,
  output [1:0]  io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_ifu_async_error_start,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [63:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [63:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_13_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_14_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_15_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_16_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_17_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_18_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_19_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_20_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_20_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_21_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_21_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_22_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_22_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_23_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_23_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_24_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_24_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_25_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_25_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_26_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_26_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_27_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_27_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_28_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_28_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_29_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_29_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_30_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_30_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_31_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_31_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_32_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_32_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_33_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_33_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_35_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_35_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_36_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_36_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_37_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_37_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_38_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_38_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_39_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_39_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_40_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_40_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_41_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_41_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_42_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_42_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_43_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_43_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_44_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_44_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_45_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_45_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_46_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_46_io_en; // @[lib.scala 343:22]
  reg  flush_final_f; // @[Reg.scala 27:20]
  wire  _T = io_exu_flush_final ^ flush_final_f; // @[lib.scala 475:21]
  wire  _T_1 = |_T; // @[lib.scala 475:29]
  reg  ifc_fetch_req_f_raw; // @[Reg.scala 27:20]
  wire  _T_339 = ~io_exu_flush_final; // @[ifu_mem_ctl.scala 225:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_339; // @[ifu_mem_ctl.scala 225:42]
  wire  _T_3 = io_ifc_fetch_req_bf_raw | ifc_fetch_req_f; // @[ifu_mem_ctl.scala 86:53]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[ifu_mem_ctl.scala 155:30]
  wire  _T_4 = _T_3 | miss_pending; // @[ifu_mem_ctl.scala 86:71]
  wire  _T_5 = _T_4 | io_exu_flush_final; // @[ifu_mem_ctl.scala 86:86]
  reg  scnd_miss_req_q; // @[Reg.scala 27:20]
  wire  scnd_miss_req = scnd_miss_req_q & _T_339; // @[ifu_mem_ctl.scala 458:36]
  wire  fetch_bf_f_c1_clken = _T_5 | scnd_miss_req; // @[ifu_mem_ctl.scala 86:107]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[ifu_mem_ctl.scala 87:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[Reg.scala 27:20]
  wire [4:0] _GEN_515 = {{1'd0}, ic_fetch_val_int_f}; // @[ifu_mem_ctl.scala 561:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_515 << ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 561:53]
  wire  _T_3199 = |ic_fetch_val_shift_right[3:2]; // @[ifu_mem_ctl.scala 563:91]
  wire  _T_3201 = _T_3199 & _T_339; // @[ifu_mem_ctl.scala 563:95]
  reg  ifc_iccm_access_f; // @[Reg.scala 27:20]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[ifu_mem_ctl.scala 177:46]
  wire  _T_3202 = _T_3201 & fetch_req_iccm_f; // @[ifu_mem_ctl.scala 563:117]
  reg  iccm_dma_rvalid_in; // @[Reg.scala 27:20]
  wire  _T_3203 = _T_3202 | iccm_dma_rvalid_in; // @[ifu_mem_ctl.scala 563:137]
  wire  _T_3204 = ~io_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[ifu_mem_ctl.scala 563:161]
  wire  _T_3205 = _T_3203 & _T_3204; // @[ifu_mem_ctl.scala 563:159]
  wire  _T_3191 = |ic_fetch_val_shift_right[1:0]; // @[ifu_mem_ctl.scala 563:91]
  wire  _T_3193 = _T_3191 & _T_339; // @[ifu_mem_ctl.scala 563:95]
  wire  _T_3194 = _T_3193 & fetch_req_iccm_f; // @[ifu_mem_ctl.scala 563:117]
  wire  _T_3195 = _T_3194 | iccm_dma_rvalid_in; // @[ifu_mem_ctl.scala 563:137]
  wire  _T_3197 = _T_3195 & _T_3204; // @[ifu_mem_ctl.scala 563:159]
  wire [1:0] iccm_ecc_word_enable = {_T_3205,_T_3197}; // @[Cat.scala 29:58]
  wire  _T_3690 = ^io_iccm_rd_data_ecc[70:39]; // @[lib.scala 193:30]
  wire  _T_3691 = ^io_iccm_rd_data_ecc[77:71]; // @[lib.scala 193:44]
  wire  _T_3692 = _T_3690 ^ _T_3691; // @[lib.scala 193:35]
  wire [5:0] _T_3700 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[lib.scala 193:76]
  wire  _T_3701 = ^_T_3700; // @[lib.scala 193:83]
  wire  _T_3702 = io_iccm_rd_data_ecc[76] ^ _T_3701; // @[lib.scala 193:71]
  wire [6:0] _T_3709 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[lib.scala 193:103]
  wire [14:0] _T_3717 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3709}; // @[lib.scala 193:103]
  wire  _T_3718 = ^_T_3717; // @[lib.scala 193:110]
  wire  _T_3719 = io_iccm_rd_data_ecc[75] ^ _T_3718; // @[lib.scala 193:98]
  wire [6:0] _T_3726 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[lib.scala 193:130]
  wire [14:0] _T_3734 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3726}; // @[lib.scala 193:130]
  wire  _T_3735 = ^_T_3734; // @[lib.scala 193:137]
  wire  _T_3736 = io_iccm_rd_data_ecc[74] ^ _T_3735; // @[lib.scala 193:125]
  wire [8:0] _T_3745 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[lib.scala 193:157]
  wire [17:0] _T_3754 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3745}; // @[lib.scala 193:157]
  wire  _T_3755 = ^_T_3754; // @[lib.scala 193:164]
  wire  _T_3756 = io_iccm_rd_data_ecc[73] ^ _T_3755; // @[lib.scala 193:152]
  wire [8:0] _T_3765 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[lib.scala 193:184]
  wire [17:0] _T_3774 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3765}; // @[lib.scala 193:184]
  wire  _T_3775 = ^_T_3774; // @[lib.scala 193:191]
  wire  _T_3776 = io_iccm_rd_data_ecc[72] ^ _T_3775; // @[lib.scala 193:179]
  wire [8:0] _T_3785 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[lib.scala 193:211]
  wire [17:0] _T_3794 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3785}; // @[lib.scala 193:211]
  wire  _T_3795 = ^_T_3794; // @[lib.scala 193:218]
  wire  _T_3796 = io_iccm_rd_data_ecc[71] ^ _T_3795; // @[lib.scala 193:206]
  wire [6:0] _T_3802 = {_T_3692,_T_3702,_T_3719,_T_3736,_T_3756,_T_3776,_T_3796}; // @[Cat.scala 29:58]
  wire  _T_3803 = _T_3802 != 7'h0; // @[lib.scala 194:44]
  wire  _T_3804 = iccm_ecc_word_enable[1] & _T_3803; // @[lib.scala 194:32]
  wire  _T_3806 = _T_3804 & _T_3802[6]; // @[lib.scala 194:53]
  wire  _T_3305 = ^io_iccm_rd_data_ecc[31:0]; // @[lib.scala 193:30]
  wire  _T_3306 = ^io_iccm_rd_data_ecc[38:32]; // @[lib.scala 193:44]
  wire  _T_3307 = _T_3305 ^ _T_3306; // @[lib.scala 193:35]
  wire [5:0] _T_3315 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[lib.scala 193:76]
  wire  _T_3316 = ^_T_3315; // @[lib.scala 193:83]
  wire  _T_3317 = io_iccm_rd_data_ecc[37] ^ _T_3316; // @[lib.scala 193:71]
  wire [6:0] _T_3324 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[lib.scala 193:103]
  wire [14:0] _T_3332 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3324}; // @[lib.scala 193:103]
  wire  _T_3333 = ^_T_3332; // @[lib.scala 193:110]
  wire  _T_3334 = io_iccm_rd_data_ecc[36] ^ _T_3333; // @[lib.scala 193:98]
  wire [6:0] _T_3341 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[lib.scala 193:130]
  wire [14:0] _T_3349 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3341}; // @[lib.scala 193:130]
  wire  _T_3350 = ^_T_3349; // @[lib.scala 193:137]
  wire  _T_3351 = io_iccm_rd_data_ecc[35] ^ _T_3350; // @[lib.scala 193:125]
  wire [8:0] _T_3360 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[lib.scala 193:157]
  wire [17:0] _T_3369 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3360}; // @[lib.scala 193:157]
  wire  _T_3370 = ^_T_3369; // @[lib.scala 193:164]
  wire  _T_3371 = io_iccm_rd_data_ecc[34] ^ _T_3370; // @[lib.scala 193:152]
  wire [8:0] _T_3380 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[lib.scala 193:184]
  wire [17:0] _T_3389 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3380}; // @[lib.scala 193:184]
  wire  _T_3390 = ^_T_3389; // @[lib.scala 193:191]
  wire  _T_3391 = io_iccm_rd_data_ecc[33] ^ _T_3390; // @[lib.scala 193:179]
  wire [8:0] _T_3400 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[lib.scala 193:211]
  wire [17:0] _T_3409 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3400}; // @[lib.scala 193:211]
  wire  _T_3410 = ^_T_3409; // @[lib.scala 193:218]
  wire  _T_3411 = io_iccm_rd_data_ecc[32] ^ _T_3410; // @[lib.scala 193:206]
  wire [6:0] _T_3417 = {_T_3307,_T_3317,_T_3334,_T_3351,_T_3371,_T_3391,_T_3411}; // @[Cat.scala 29:58]
  wire  _T_3418 = _T_3417 != 7'h0; // @[lib.scala 194:44]
  wire  _T_3419 = iccm_ecc_word_enable[0] & _T_3418; // @[lib.scala 194:32]
  wire  _T_3421 = _T_3419 & _T_3417[6]; // @[lib.scala 194:53]
  wire [1:0] iccm_single_ecc_error = {_T_3806,_T_3421}; // @[Cat.scala 29:58]
  wire  _T_6 = |iccm_single_ecc_error; // @[ifu_mem_ctl.scala 91:52]
  reg  dma_iccm_req_f; // @[Reg.scala 27:20]
  wire  _T_9 = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err | io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu_mem_ctl.scala 92:74]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_10 = perr_state == 3'h4; // @[ifu_mem_ctl.scala 93:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[ifu_mem_ctl.scala 383:34]
  wire  _T_11 = iccm_correct_ecc | _T_10; // @[ifu_mem_ctl.scala 93:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_12 = err_stop_state == 2'h3; // @[ifu_mem_ctl.scala 93:90]
  wire  _T_13 = _T_11 | _T_12; // @[ifu_mem_ctl.scala 93:72]
  wire  _T_2547 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2552 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2572 = io_ifu_fetch_val == 2'h3; // @[ifu_mem_ctl.scala 430:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[ifu_mem_ctl.scala 297:42]
  wire  _T_2574 = io_ifu_fetch_val[0] & two_byte_instr; // @[ifu_mem_ctl.scala 430:79]
  wire  _T_2575 = _T_2572 | _T_2574; // @[ifu_mem_ctl.scala 430:56]
  wire  _T_2576 = io_exu_flush_final | io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 430:122]
  wire  _T_2577 = ~_T_2576; // @[ifu_mem_ctl.scala 430:101]
  wire  _T_2578 = _T_2575 & _T_2577; // @[ifu_mem_ctl.scala 430:99]
  wire  _T_2579 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2593 = io_ifu_fetch_val[0] & _T_339; // @[ifu_mem_ctl.scala 437:45]
  wire  _T_2594 = ~io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 437:69]
  wire  _T_2595 = _T_2593 & _T_2594; // @[ifu_mem_ctl.scala 437:67]
  wire  _T_2596 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_76 = _T_2579 ? _T_2595 : _T_2596; // @[Conditional.scala 39:67]
  wire  _GEN_80 = _T_2552 ? _T_2578 : _GEN_76; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2547 ? 1'h0 : _GEN_80; // @[Conditional.scala 40:58]
  wire  _T_14 = _T_13 | err_stop_fetch; // @[ifu_mem_ctl.scala 93:112]
  wire  _T_16 = io_ifu_axi_r_valid & io_ifu_bus_clk_en; // @[ifu_mem_ctl.scala 95:45]
  wire  _T_17 = _T_16 & io_ifu_axi_r_ready; // @[ifu_mem_ctl.scala 95:66]
  wire  _T_233 = |io_ic_rd_hit; // @[ifu_mem_ctl.scala 185:37]
  wire  _T_234 = ~_T_233; // @[ifu_mem_ctl.scala 185:23]
  reg  reset_all_tags; // @[Reg.scala 27:20]
  wire  _T_235 = _T_234 | reset_all_tags; // @[ifu_mem_ctl.scala 185:41]
  wire  _T_213 = ~ifc_iccm_access_f; // @[ifu_mem_ctl.scala 176:48]
  wire  _T_214 = ifc_fetch_req_f & _T_213; // @[ifu_mem_ctl.scala 176:46]
  reg  ifc_region_acc_fault_final_f; // @[Reg.scala 27:20]
  wire  _T_215 = ~ifc_region_acc_fault_final_f; // @[ifu_mem_ctl.scala 176:69]
  wire  fetch_req_icache_f = _T_214 & _T_215; // @[ifu_mem_ctl.scala 176:67]
  wire  _T_236 = _T_235 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 185:59]
  wire  _T_237 = ~miss_pending; // @[ifu_mem_ctl.scala 185:82]
  wire  _T_238 = _T_236 & _T_237; // @[ifu_mem_ctl.scala 185:80]
  wire  _T_239 = _T_238 | scnd_miss_req; // @[ifu_mem_ctl.scala 185:97]
  wire  ic_act_miss_f = _T_239 & _T_215; // @[ifu_mem_ctl.scala 185:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[ifu_mem_ctl.scala 488:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[ifu_mem_ctl.scala 516:41]
  reg  uncacheable_miss_ff; // @[Reg.scala 27:20]
  reg [2:0] bus_data_beat_count; // @[Reg.scala 27:20]
  wire  _T_2713 = bus_data_beat_count == 3'h1; // @[ifu_mem_ctl.scala 514:69]
  wire  _T_2714 = &bus_data_beat_count; // @[ifu_mem_ctl.scala 514:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2713 : _T_2714; // @[ifu_mem_ctl.scala 514:28]
  wire  _T_2654 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[ifu_mem_ctl.scala 493:68]
  wire  _T_2655 = ic_act_miss_f | _T_2654; // @[ifu_mem_ctl.scala 493:48]
  wire  bus_reset_data_beat_cnt = _T_2655 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 493:91]
  wire  _T_2651 = ~bus_last_data_beat; // @[ifu_mem_ctl.scala 492:50]
  wire  _T_2652 = bus_ifu_wr_en_ff & _T_2651; // @[ifu_mem_ctl.scala 492:48]
  wire  _T_2653 = ~io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 492:72]
  wire  bus_inc_data_beat_cnt = _T_2652 & _T_2653; // @[ifu_mem_ctl.scala 492:70]
  wire [2:0] _T_2659 = bus_data_beat_count + 3'h1; // @[ifu_mem_ctl.scala 496:115]
  wire [2:0] _T_2661 = bus_inc_data_beat_cnt ? _T_2659 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2656 = ~bus_inc_data_beat_cnt; // @[ifu_mem_ctl.scala 494:32]
  wire  _T_2657 = ~bus_reset_data_beat_cnt; // @[ifu_mem_ctl.scala 494:57]
  wire  bus_hold_data_beat_cnt = _T_2656 & _T_2657; // @[ifu_mem_ctl.scala 494:55]
  wire [2:0] _T_2662 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2661 | _T_2662; // @[Mux.scala 27:72]
  wire  _T_18 = &bus_new_data_beat_count; // @[ifu_mem_ctl.scala 95:114]
  wire  _T_19 = _T_17 & _T_18; // @[ifu_mem_ctl.scala 95:87]
  wire  _T_20 = ~uncacheable_miss_ff; // @[ifu_mem_ctl.scala 96:5]
  wire  _T_21 = _T_19 & _T_20; // @[ifu_mem_ctl.scala 95:120]
  wire  _T_22 = miss_state == 3'h5; // @[ifu_mem_ctl.scala 96:41]
  wire  _T_27 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_29 = ic_act_miss_f & _T_339; // @[ifu_mem_ctl.scala 102:43]
  wire [2:0] _T_31 = _T_29 ? 3'h1 : 3'h2; // @[ifu_mem_ctl.scala 102:27]
  wire  _T_34 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[ifu_mem_ctl.scala 333:45]
  wire  _T_2161 = byp_fetch_index[4:2] == 3'h0; // @[ifu_mem_ctl.scala 353:127]
  reg [7:0] ic_miss_buff_data_valid; // @[ifu_mem_ctl.scala 310:62]
  wire  _T_2192 = _T_2161 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2165 = byp_fetch_index[4:2] == 3'h1; // @[ifu_mem_ctl.scala 353:127]
  wire  _T_2193 = _T_2165 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2200 = _T_2192 | _T_2193; // @[Mux.scala 27:72]
  wire  _T_2169 = byp_fetch_index[4:2] == 3'h2; // @[ifu_mem_ctl.scala 353:127]
  wire  _T_2194 = _T_2169 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2201 = _T_2200 | _T_2194; // @[Mux.scala 27:72]
  wire  _T_2173 = byp_fetch_index[4:2] == 3'h3; // @[ifu_mem_ctl.scala 353:127]
  wire  _T_2195 = _T_2173 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2202 = _T_2201 | _T_2195; // @[Mux.scala 27:72]
  wire  _T_2177 = byp_fetch_index[4:2] == 3'h4; // @[ifu_mem_ctl.scala 353:127]
  wire  _T_2196 = _T_2177 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2203 = _T_2202 | _T_2196; // @[Mux.scala 27:72]
  wire  _T_2181 = byp_fetch_index[4:2] == 3'h5; // @[ifu_mem_ctl.scala 353:127]
  wire  _T_2197 = _T_2181 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2204 = _T_2203 | _T_2197; // @[Mux.scala 27:72]
  wire  _T_2185 = byp_fetch_index[4:2] == 3'h6; // @[ifu_mem_ctl.scala 353:127]
  wire  _T_2198 = _T_2185 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2205 = _T_2204 | _T_2198; // @[Mux.scala 27:72]
  wire  _T_2189 = byp_fetch_index[4:2] == 3'h7; // @[ifu_mem_ctl.scala 353:127]
  wire  _T_2199 = _T_2189 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2205 | _T_2199; // @[Mux.scala 27:72]
  wire  _T_2247 = ~byp_fetch_index[1]; // @[ifu_mem_ctl.scala 355:69]
  wire  _T_2248 = ic_miss_buff_data_valid_bypass_index & _T_2247; // @[ifu_mem_ctl.scala 355:67]
  wire  _T_2250 = ~byp_fetch_index[0]; // @[ifu_mem_ctl.scala 355:91]
  wire  _T_2251 = _T_2248 & _T_2250; // @[ifu_mem_ctl.scala 355:89]
  wire  _T_2256 = _T_2248 & byp_fetch_index[0]; // @[ifu_mem_ctl.scala 356:65]
  wire  _T_2257 = _T_2251 | _T_2256; // @[ifu_mem_ctl.scala 355:112]
  wire  _T_2259 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[ifu_mem_ctl.scala 357:43]
  wire  _T_2262 = _T_2259 & _T_2250; // @[ifu_mem_ctl.scala 357:65]
  wire  _T_2263 = _T_2257 | _T_2262; // @[ifu_mem_ctl.scala 356:88]
  wire  _T_2267 = _T_2259 & byp_fetch_index[0]; // @[ifu_mem_ctl.scala 358:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[ifu_mem_ctl.scala 336:75]
  wire  _T_2207 = byp_fetch_index_inc == 3'h0; // @[ifu_mem_ctl.scala 354:110]
  wire  _T_2231 = _T_2207 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2210 = byp_fetch_index_inc == 3'h1; // @[ifu_mem_ctl.scala 354:110]
  wire  _T_2232 = _T_2210 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2239 = _T_2231 | _T_2232; // @[Mux.scala 27:72]
  wire  _T_2213 = byp_fetch_index_inc == 3'h2; // @[ifu_mem_ctl.scala 354:110]
  wire  _T_2233 = _T_2213 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2240 = _T_2239 | _T_2233; // @[Mux.scala 27:72]
  wire  _T_2216 = byp_fetch_index_inc == 3'h3; // @[ifu_mem_ctl.scala 354:110]
  wire  _T_2234 = _T_2216 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2241 = _T_2240 | _T_2234; // @[Mux.scala 27:72]
  wire  _T_2219 = byp_fetch_index_inc == 3'h4; // @[ifu_mem_ctl.scala 354:110]
  wire  _T_2235 = _T_2219 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2242 = _T_2241 | _T_2235; // @[Mux.scala 27:72]
  wire  _T_2222 = byp_fetch_index_inc == 3'h5; // @[ifu_mem_ctl.scala 354:110]
  wire  _T_2236 = _T_2222 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2243 = _T_2242 | _T_2236; // @[Mux.scala 27:72]
  wire  _T_2225 = byp_fetch_index_inc == 3'h6; // @[ifu_mem_ctl.scala 354:110]
  wire  _T_2237 = _T_2225 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2244 = _T_2243 | _T_2237; // @[Mux.scala 27:72]
  wire  _T_2228 = byp_fetch_index_inc == 3'h7; // @[ifu_mem_ctl.scala 354:110]
  wire  _T_2238 = _T_2228 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2244 | _T_2238; // @[Mux.scala 27:72]
  wire  _T_2268 = _T_2267 & ic_miss_buff_data_valid_inc_bypass_index; // @[ifu_mem_ctl.scala 358:87]
  wire  _T_2269 = _T_2263 | _T_2268; // @[ifu_mem_ctl.scala 357:88]
  wire  _T_2273 = ic_miss_buff_data_valid_bypass_index & _T_2189; // @[ifu_mem_ctl.scala 359:43]
  wire  miss_buff_hit_unq_f = _T_2269 | _T_2273; // @[ifu_mem_ctl.scala 358:131]
  wire  _T_2289 = miss_state == 3'h4; // @[ifu_mem_ctl.scala 364:55]
  wire  _T_2290 = miss_state == 3'h1; // @[ifu_mem_ctl.scala 364:87]
  wire  _T_2291 = _T_2289 | _T_2290; // @[ifu_mem_ctl.scala 364:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2291; // @[ifu_mem_ctl.scala 364:41]
  wire  _T_2274 = miss_state == 3'h6; // @[ifu_mem_ctl.scala 361:30]
  reg [30:0] imb_ff; // @[Reg.scala 27:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[ifu_mem_ctl.scala 352:48]
  wire  _T_2275 = ~miss_wrap_f; // @[ifu_mem_ctl.scala 361:68]
  wire  _T_2276 = miss_buff_hit_unq_f & _T_2275; // @[ifu_mem_ctl.scala 361:66]
  wire  stream_hit_f = _T_2274 & _T_2276; // @[ifu_mem_ctl.scala 361:43]
  wire  _T_221 = crit_byp_hit_f | stream_hit_f; // @[ifu_mem_ctl.scala 180:35]
  wire  _T_222 = _T_221 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 180:52]
  wire  ic_byp_hit_f = _T_222 & miss_pending; // @[ifu_mem_ctl.scala 180:73]
  reg  last_data_recieved_ff; // @[Reg.scala 27:20]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[ifu_mem_ctl.scala 526:35]
  wire  _T_35 = bus_ifu_wr_en_ff & last_beat; // @[ifu_mem_ctl.scala 106:126]
  wire  _T_36 = last_data_recieved_ff | _T_35; // @[ifu_mem_ctl.scala 106:106]
  wire  _T_37 = ic_byp_hit_f & _T_36; // @[ifu_mem_ctl.scala 106:80]
  wire  _T_38 = _T_37 & uncacheable_miss_ff; // @[ifu_mem_ctl.scala 106:140]
  wire  _T_39 = io_dec_mem_ctrl_dec_tlu_force_halt | _T_38; // @[ifu_mem_ctl.scala 106:64]
  wire  _T_41 = ~last_data_recieved_ff; // @[ifu_mem_ctl.scala 107:30]
  wire  _T_42 = ic_byp_hit_f & _T_41; // @[ifu_mem_ctl.scala 107:27]
  wire  _T_43 = _T_42 & uncacheable_miss_ff; // @[ifu_mem_ctl.scala 107:53]
  wire  _T_45 = ~ic_byp_hit_f; // @[ifu_mem_ctl.scala 108:16]
  wire  _T_47 = _T_45 & _T_339; // @[ifu_mem_ctl.scala 108:30]
  wire  _T_49 = _T_47 & _T_35; // @[ifu_mem_ctl.scala 108:52]
  wire  _T_50 = _T_49 & uncacheable_miss_ff; // @[ifu_mem_ctl.scala 108:85]
  wire  _T_54 = _T_35 & _T_20; // @[ifu_mem_ctl.scala 109:49]
  wire  _T_57 = ic_byp_hit_f & _T_339; // @[ifu_mem_ctl.scala 110:33]
  wire  _T_59 = ~_T_35; // @[ifu_mem_ctl.scala 110:57]
  wire  _T_60 = _T_57 & _T_59; // @[ifu_mem_ctl.scala 110:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[ifu_mem_ctl.scala 98:52]
  wire  _T_61 = ~ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 110:91]
  wire  _T_62 = _T_60 & _T_61; // @[ifu_mem_ctl.scala 110:89]
  wire  _T_64 = _T_62 & _T_20; // @[ifu_mem_ctl.scala 110:113]
  wire  _T_67 = bus_ifu_wr_en_ff & _T_339; // @[ifu_mem_ctl.scala 111:39]
  wire  _T_70 = _T_67 & _T_59; // @[ifu_mem_ctl.scala 111:61]
  wire  _T_72 = _T_70 & _T_61; // @[ifu_mem_ctl.scala 111:95]
  wire  _T_74 = _T_72 & _T_20; // @[ifu_mem_ctl.scala 111:119]
  wire  _T_82 = _T_49 & _T_20; // @[ifu_mem_ctl.scala 112:102]
  wire  _T_84 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 113:46]
  wire  _T_87 = _T_84 & _T_59; // @[ifu_mem_ctl.scala 113:70]
  wire [2:0] _T_89 = _T_87 ? 3'h2 : 3'h0; // @[ifu_mem_ctl.scala 113:24]
  wire [2:0] _T_90 = _T_82 ? 3'h0 : _T_89; // @[ifu_mem_ctl.scala 112:22]
  wire [2:0] _T_91 = _T_74 ? 3'h6 : _T_90; // @[ifu_mem_ctl.scala 111:20]
  wire [2:0] _T_92 = _T_64 ? 3'h6 : _T_91; // @[ifu_mem_ctl.scala 110:18]
  wire [2:0] _T_93 = _T_54 ? 3'h0 : _T_92; // @[ifu_mem_ctl.scala 109:16]
  wire [2:0] _T_94 = _T_50 ? 3'h4 : _T_93; // @[ifu_mem_ctl.scala 108:14]
  wire [2:0] _T_95 = _T_43 ? 3'h3 : _T_94; // @[ifu_mem_ctl.scala 107:12]
  wire [2:0] _T_96 = _T_39 ? 3'h0 : _T_95; // @[ifu_mem_ctl.scala 106:27]
  wire  _T_105 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_109 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2286 = byp_fetch_index[4:1] == 4'hf; // @[ifu_mem_ctl.scala 363:60]
  wire  _T_2287 = _T_2286 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 363:94]
  wire  stream_eol_f = _T_2287 & stream_hit_f; // @[ifu_mem_ctl.scala 363:112]
  wire  _T_111 = _T_84 | stream_eol_f; // @[ifu_mem_ctl.scala 121:72]
  wire  _T_114 = _T_111 & _T_59; // @[ifu_mem_ctl.scala 121:87]
  wire  _T_116 = _T_114 & _T_2653; // @[ifu_mem_ctl.scala 121:122]
  wire [2:0] _T_118 = _T_116 ? 3'h2 : 3'h0; // @[ifu_mem_ctl.scala 121:27]
  wire  _T_124 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_127 = io_exu_flush_final & _T_59; // @[ifu_mem_ctl.scala 125:48]
  wire  _T_129 = _T_127 & _T_2653; // @[ifu_mem_ctl.scala 125:82]
  wire [2:0] _T_131 = _T_129 ? 3'h2 : 3'h0; // @[ifu_mem_ctl.scala 125:27]
  wire  _T_135 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_242 = io_ic_rd_hit == 2'h0; // @[ifu_mem_ctl.scala 186:28]
  wire  _T_243 = _T_242 | reset_all_tags; // @[ifu_mem_ctl.scala 186:42]
  wire  _T_244 = _T_243 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 186:60]
  wire  _T_245 = miss_state == 3'h2; // @[ifu_mem_ctl.scala 186:94]
  wire  _T_246 = _T_244 & _T_245; // @[ifu_mem_ctl.scala 186:81]
  wire  _T_249 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[ifu_mem_ctl.scala 187:39]
  wire  _T_250 = _T_246 & _T_249; // @[ifu_mem_ctl.scala 186:111]
  wire  _T_252 = _T_250 & _T_20; // @[ifu_mem_ctl.scala 187:91]
  reg  sel_mb_addr_ff; // @[Reg.scala 27:20]
  wire  _T_253 = ~sel_mb_addr_ff; // @[ifu_mem_ctl.scala 187:116]
  wire  _T_254 = _T_252 & _T_253; // @[ifu_mem_ctl.scala 187:114]
  wire  ic_miss_under_miss_f = _T_254 & _T_215; // @[ifu_mem_ctl.scala 187:132]
  wire  _T_138 = ic_miss_under_miss_f & _T_59; // @[ifu_mem_ctl.scala 129:50]
  wire  _T_140 = _T_138 & _T_2653; // @[ifu_mem_ctl.scala 129:84]
  wire  _T_262 = _T_236 & _T_245; // @[ifu_mem_ctl.scala 188:85]
  wire  _T_265 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[ifu_mem_ctl.scala 189:39]
  wire  _T_266 = _T_265 | uncacheable_miss_ff; // @[ifu_mem_ctl.scala 189:91]
  wire  ic_ignore_2nd_miss_f = _T_262 & _T_266; // @[ifu_mem_ctl.scala 188:117]
  wire  _T_144 = ic_ignore_2nd_miss_f & _T_59; // @[ifu_mem_ctl.scala 130:35]
  wire  _T_146 = _T_144 & _T_2653; // @[ifu_mem_ctl.scala 130:69]
  wire [2:0] _T_148 = _T_146 ? 3'h7 : 3'h0; // @[ifu_mem_ctl.scala 130:12]
  wire [2:0] _T_149 = _T_140 ? 3'h5 : _T_148; // @[ifu_mem_ctl.scala 129:27]
  wire  _T_154 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_157 = _T_35 ? 3'h0 : 3'h2; // @[ifu_mem_ctl.scala 135:12]
  wire [2:0] _T_158 = io_exu_flush_final ? _T_157 : 3'h1; // @[ifu_mem_ctl.scala 134:75]
  wire [2:0] _T_159 = io_dec_mem_ctrl_dec_tlu_force_halt ? 3'h0 : _T_158; // @[ifu_mem_ctl.scala 134:27]
  wire  _T_163 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_167 = io_exu_flush_final ? _T_157 : 3'h0; // @[ifu_mem_ctl.scala 139:75]
  wire [2:0] _T_168 = io_dec_mem_ctrl_dec_tlu_force_halt ? 3'h0 : _T_167; // @[ifu_mem_ctl.scala 139:27]
  wire [2:0] _GEN_1 = _T_163 ? _T_168 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_3 = _T_154 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_5 = _T_135 ? _T_149 : _GEN_3; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_7 = _T_124 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_9 = _T_109 ? _T_118 : _GEN_7; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_11 = _T_105 ? 3'h0 : _GEN_9; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_13 = _T_34 ? _T_96 : _GEN_11; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_27 ? _T_31 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_23 = miss_nxtstate == 3'h5; // @[ifu_mem_ctl.scala 96:73]
  wire  _T_24 = _T_22 | _T_23; // @[ifu_mem_ctl.scala 96:57]
  wire  _T_25 = _T_21 & _T_24; // @[ifu_mem_ctl.scala 96:26]
  wire  scnd_miss_req_in = _T_25 & _T_339; // @[ifu_mem_ctl.scala 96:91]
  wire  _T_33 = ic_act_miss_f & _T_2653; // @[ifu_mem_ctl.scala 103:38]
  wire  _T_97 = io_dec_mem_ctrl_dec_tlu_force_halt | io_exu_flush_final; // @[ifu_mem_ctl.scala 114:59]
  wire  _T_98 = _T_97 | ic_byp_hit_f; // @[ifu_mem_ctl.scala 114:80]
  wire  _T_99 = _T_98 | ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 114:95]
  wire  _T_101 = _T_99 | _T_35; // @[ifu_mem_ctl.scala 114:118]
  wire  _T_103 = bus_ifu_wr_en_ff & _T_20; // @[ifu_mem_ctl.scala 114:171]
  wire  _T_104 = _T_101 | _T_103; // @[ifu_mem_ctl.scala 114:151]
  wire  _T_106 = io_exu_flush_final | flush_final_f; // @[ifu_mem_ctl.scala 118:43]
  wire  _T_107 = _T_106 | ic_byp_hit_f; // @[ifu_mem_ctl.scala 118:59]
  wire  _T_108 = _T_107 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 118:74]
  wire  _T_122 = _T_111 | _T_35; // @[ifu_mem_ctl.scala 122:84]
  wire  _T_123 = _T_122 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 122:118]
  wire  _T_133 = io_exu_flush_final | _T_35; // @[ifu_mem_ctl.scala 126:43]
  wire  _T_134 = _T_133 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 126:76]
  wire  _T_151 = _T_35 | ic_miss_under_miss_f; // @[ifu_mem_ctl.scala 131:55]
  wire  _T_152 = _T_151 | ic_ignore_2nd_miss_f; // @[ifu_mem_ctl.scala 131:78]
  wire  _T_153 = _T_152 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 131:101]
  wire  _T_161 = _T_35 | io_exu_flush_final; // @[ifu_mem_ctl.scala 136:55]
  wire  _T_162 = _T_161 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 136:76]
  wire  _GEN_2 = _T_163 & _T_162; // @[Conditional.scala 39:67]
  wire  _GEN_4 = _T_154 ? _T_162 : _GEN_2; // @[Conditional.scala 39:67]
  wire  _GEN_6 = _T_135 ? _T_153 : _GEN_4; // @[Conditional.scala 39:67]
  wire  _GEN_8 = _T_124 ? _T_134 : _GEN_6; // @[Conditional.scala 39:67]
  wire  _GEN_10 = _T_109 ? _T_123 : _GEN_8; // @[Conditional.scala 39:67]
  wire  _GEN_12 = _T_105 ? _T_108 : _GEN_10; // @[Conditional.scala 39:67]
  wire  _GEN_14 = _T_34 ? _T_104 : _GEN_12; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_27 ? _T_33 : _GEN_14; // @[Conditional.scala 40:58]
  wire  _T_177 = ~flush_final_f; // @[ifu_mem_ctl.scala 156:95]
  wire  _T_178 = _T_2289 & _T_177; // @[ifu_mem_ctl.scala 156:93]
  wire  crit_wd_byp_ok_ff = _T_2290 | _T_178; // @[ifu_mem_ctl.scala 156:58]
  wire  _T_181 = miss_pending & _T_59; // @[ifu_mem_ctl.scala 157:36]
  wire  _T_183 = _T_2289 & io_exu_flush_final; // @[ifu_mem_ctl.scala 157:106]
  wire  _T_184 = ~_T_183; // @[ifu_mem_ctl.scala 157:72]
  wire  _T_185 = _T_181 & _T_184; // @[ifu_mem_ctl.scala 157:70]
  wire  _T_187 = _T_2289 & crit_byp_hit_f; // @[ifu_mem_ctl.scala 158:39]
  wire  _T_188 = ~_T_187; // @[ifu_mem_ctl.scala 158:5]
  wire  _T_189 = _T_185 & _T_188; // @[ifu_mem_ctl.scala 157:128]
  wire  _T_190 = _T_189 | ic_act_miss_f; // @[ifu_mem_ctl.scala 158:59]
  wire  _T_191 = miss_nxtstate == 3'h4; // @[ifu_mem_ctl.scala 159:36]
  wire  _T_192 = miss_pending & _T_191; // @[ifu_mem_ctl.scala 159:19]
  wire  sel_hold_imb = _T_190 | _T_192; // @[ifu_mem_ctl.scala 158:75]
  wire  _T_194 = _T_22 | ic_miss_under_miss_f; // @[ifu_mem_ctl.scala 161:57]
  wire  sel_hold_imb_scnd = _T_194 & _T_177; // @[ifu_mem_ctl.scala 161:81]
  reg  way_status_mb_scnd_ff; // @[Reg.scala 27:20]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[Reg.scala 27:20]
  wire  _T_4900 = ifu_ic_rw_int_addr_ff == 7'h0; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire  _T_5028 = _T_4900 & way_status_out_0; // @[Mux.scala 27:72]
  wire  _T_4901 = ifu_ic_rw_int_addr_ff == 7'h1; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire  _T_5029 = _T_4901 & way_status_out_1; // @[Mux.scala 27:72]
  wire  _T_5156 = _T_5028 | _T_5029; // @[Mux.scala 27:72]
  wire  _T_4902 = ifu_ic_rw_int_addr_ff == 7'h2; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire  _T_5030 = _T_4902 & way_status_out_2; // @[Mux.scala 27:72]
  wire  _T_5157 = _T_5156 | _T_5030; // @[Mux.scala 27:72]
  wire  _T_4903 = ifu_ic_rw_int_addr_ff == 7'h3; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire  _T_5031 = _T_4903 & way_status_out_3; // @[Mux.scala 27:72]
  wire  _T_5158 = _T_5157 | _T_5031; // @[Mux.scala 27:72]
  wire  _T_4904 = ifu_ic_rw_int_addr_ff == 7'h4; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire  _T_5032 = _T_4904 & way_status_out_4; // @[Mux.scala 27:72]
  wire  _T_5159 = _T_5158 | _T_5032; // @[Mux.scala 27:72]
  wire  _T_4905 = ifu_ic_rw_int_addr_ff == 7'h5; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire  _T_5033 = _T_4905 & way_status_out_5; // @[Mux.scala 27:72]
  wire  _T_5160 = _T_5159 | _T_5033; // @[Mux.scala 27:72]
  wire  _T_4906 = ifu_ic_rw_int_addr_ff == 7'h6; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire  _T_5034 = _T_4906 & way_status_out_6; // @[Mux.scala 27:72]
  wire  _T_5161 = _T_5160 | _T_5034; // @[Mux.scala 27:72]
  wire  _T_4907 = ifu_ic_rw_int_addr_ff == 7'h7; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire  _T_5035 = _T_4907 & way_status_out_7; // @[Mux.scala 27:72]
  wire  _T_5162 = _T_5161 | _T_5035; // @[Mux.scala 27:72]
  wire  _T_4908 = ifu_ic_rw_int_addr_ff == 7'h8; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire  _T_5036 = _T_4908 & way_status_out_8; // @[Mux.scala 27:72]
  wire  _T_5163 = _T_5162 | _T_5036; // @[Mux.scala 27:72]
  wire  _T_4909 = ifu_ic_rw_int_addr_ff == 7'h9; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire  _T_5037 = _T_4909 & way_status_out_9; // @[Mux.scala 27:72]
  wire  _T_5164 = _T_5163 | _T_5037; // @[Mux.scala 27:72]
  wire  _T_4910 = ifu_ic_rw_int_addr_ff == 7'ha; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire  _T_5038 = _T_4910 & way_status_out_10; // @[Mux.scala 27:72]
  wire  _T_5165 = _T_5164 | _T_5038; // @[Mux.scala 27:72]
  wire  _T_4911 = ifu_ic_rw_int_addr_ff == 7'hb; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire  _T_5039 = _T_4911 & way_status_out_11; // @[Mux.scala 27:72]
  wire  _T_5166 = _T_5165 | _T_5039; // @[Mux.scala 27:72]
  wire  _T_4912 = ifu_ic_rw_int_addr_ff == 7'hc; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire  _T_5040 = _T_4912 & way_status_out_12; // @[Mux.scala 27:72]
  wire  _T_5167 = _T_5166 | _T_5040; // @[Mux.scala 27:72]
  wire  _T_4913 = ifu_ic_rw_int_addr_ff == 7'hd; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire  _T_5041 = _T_4913 & way_status_out_13; // @[Mux.scala 27:72]
  wire  _T_5168 = _T_5167 | _T_5041; // @[Mux.scala 27:72]
  wire  _T_4914 = ifu_ic_rw_int_addr_ff == 7'he; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire  _T_5042 = _T_4914 & way_status_out_14; // @[Mux.scala 27:72]
  wire  _T_5169 = _T_5168 | _T_5042; // @[Mux.scala 27:72]
  wire  _T_4915 = ifu_ic_rw_int_addr_ff == 7'hf; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire  _T_5043 = _T_4915 & way_status_out_15; // @[Mux.scala 27:72]
  wire  _T_5170 = _T_5169 | _T_5043; // @[Mux.scala 27:72]
  wire  _T_4916 = ifu_ic_rw_int_addr_ff == 7'h10; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire  _T_5044 = _T_4916 & way_status_out_16; // @[Mux.scala 27:72]
  wire  _T_5171 = _T_5170 | _T_5044; // @[Mux.scala 27:72]
  wire  _T_4917 = ifu_ic_rw_int_addr_ff == 7'h11; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire  _T_5045 = _T_4917 & way_status_out_17; // @[Mux.scala 27:72]
  wire  _T_5172 = _T_5171 | _T_5045; // @[Mux.scala 27:72]
  wire  _T_4918 = ifu_ic_rw_int_addr_ff == 7'h12; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire  _T_5046 = _T_4918 & way_status_out_18; // @[Mux.scala 27:72]
  wire  _T_5173 = _T_5172 | _T_5046; // @[Mux.scala 27:72]
  wire  _T_4919 = ifu_ic_rw_int_addr_ff == 7'h13; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire  _T_5047 = _T_4919 & way_status_out_19; // @[Mux.scala 27:72]
  wire  _T_5174 = _T_5173 | _T_5047; // @[Mux.scala 27:72]
  wire  _T_4920 = ifu_ic_rw_int_addr_ff == 7'h14; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire  _T_5048 = _T_4920 & way_status_out_20; // @[Mux.scala 27:72]
  wire  _T_5175 = _T_5174 | _T_5048; // @[Mux.scala 27:72]
  wire  _T_4921 = ifu_ic_rw_int_addr_ff == 7'h15; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire  _T_5049 = _T_4921 & way_status_out_21; // @[Mux.scala 27:72]
  wire  _T_5176 = _T_5175 | _T_5049; // @[Mux.scala 27:72]
  wire  _T_4922 = ifu_ic_rw_int_addr_ff == 7'h16; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire  _T_5050 = _T_4922 & way_status_out_22; // @[Mux.scala 27:72]
  wire  _T_5177 = _T_5176 | _T_5050; // @[Mux.scala 27:72]
  wire  _T_4923 = ifu_ic_rw_int_addr_ff == 7'h17; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire  _T_5051 = _T_4923 & way_status_out_23; // @[Mux.scala 27:72]
  wire  _T_5178 = _T_5177 | _T_5051; // @[Mux.scala 27:72]
  wire  _T_4924 = ifu_ic_rw_int_addr_ff == 7'h18; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire  _T_5052 = _T_4924 & way_status_out_24; // @[Mux.scala 27:72]
  wire  _T_5179 = _T_5178 | _T_5052; // @[Mux.scala 27:72]
  wire  _T_4925 = ifu_ic_rw_int_addr_ff == 7'h19; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire  _T_5053 = _T_4925 & way_status_out_25; // @[Mux.scala 27:72]
  wire  _T_5180 = _T_5179 | _T_5053; // @[Mux.scala 27:72]
  wire  _T_4926 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire  _T_5054 = _T_4926 & way_status_out_26; // @[Mux.scala 27:72]
  wire  _T_5181 = _T_5180 | _T_5054; // @[Mux.scala 27:72]
  wire  _T_4927 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire  _T_5055 = _T_4927 & way_status_out_27; // @[Mux.scala 27:72]
  wire  _T_5182 = _T_5181 | _T_5055; // @[Mux.scala 27:72]
  wire  _T_4928 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire  _T_5056 = _T_4928 & way_status_out_28; // @[Mux.scala 27:72]
  wire  _T_5183 = _T_5182 | _T_5056; // @[Mux.scala 27:72]
  wire  _T_4929 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire  _T_5057 = _T_4929 & way_status_out_29; // @[Mux.scala 27:72]
  wire  _T_5184 = _T_5183 | _T_5057; // @[Mux.scala 27:72]
  wire  _T_4930 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire  _T_5058 = _T_4930 & way_status_out_30; // @[Mux.scala 27:72]
  wire  _T_5185 = _T_5184 | _T_5058; // @[Mux.scala 27:72]
  wire  _T_4931 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire  _T_5059 = _T_4931 & way_status_out_31; // @[Mux.scala 27:72]
  wire  _T_5186 = _T_5185 | _T_5059; // @[Mux.scala 27:72]
  wire  _T_4932 = ifu_ic_rw_int_addr_ff == 7'h20; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire  _T_5060 = _T_4932 & way_status_out_32; // @[Mux.scala 27:72]
  wire  _T_5187 = _T_5186 | _T_5060; // @[Mux.scala 27:72]
  wire  _T_4933 = ifu_ic_rw_int_addr_ff == 7'h21; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire  _T_5061 = _T_4933 & way_status_out_33; // @[Mux.scala 27:72]
  wire  _T_5188 = _T_5187 | _T_5061; // @[Mux.scala 27:72]
  wire  _T_4934 = ifu_ic_rw_int_addr_ff == 7'h22; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire  _T_5062 = _T_4934 & way_status_out_34; // @[Mux.scala 27:72]
  wire  _T_5189 = _T_5188 | _T_5062; // @[Mux.scala 27:72]
  wire  _T_4935 = ifu_ic_rw_int_addr_ff == 7'h23; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire  _T_5063 = _T_4935 & way_status_out_35; // @[Mux.scala 27:72]
  wire  _T_5190 = _T_5189 | _T_5063; // @[Mux.scala 27:72]
  wire  _T_4936 = ifu_ic_rw_int_addr_ff == 7'h24; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire  _T_5064 = _T_4936 & way_status_out_36; // @[Mux.scala 27:72]
  wire  _T_5191 = _T_5190 | _T_5064; // @[Mux.scala 27:72]
  wire  _T_4937 = ifu_ic_rw_int_addr_ff == 7'h25; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire  _T_5065 = _T_4937 & way_status_out_37; // @[Mux.scala 27:72]
  wire  _T_5192 = _T_5191 | _T_5065; // @[Mux.scala 27:72]
  wire  _T_4938 = ifu_ic_rw_int_addr_ff == 7'h26; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire  _T_5066 = _T_4938 & way_status_out_38; // @[Mux.scala 27:72]
  wire  _T_5193 = _T_5192 | _T_5066; // @[Mux.scala 27:72]
  wire  _T_4939 = ifu_ic_rw_int_addr_ff == 7'h27; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire  _T_5067 = _T_4939 & way_status_out_39; // @[Mux.scala 27:72]
  wire  _T_5194 = _T_5193 | _T_5067; // @[Mux.scala 27:72]
  wire  _T_4940 = ifu_ic_rw_int_addr_ff == 7'h28; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire  _T_5068 = _T_4940 & way_status_out_40; // @[Mux.scala 27:72]
  wire  _T_5195 = _T_5194 | _T_5068; // @[Mux.scala 27:72]
  wire  _T_4941 = ifu_ic_rw_int_addr_ff == 7'h29; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire  _T_5069 = _T_4941 & way_status_out_41; // @[Mux.scala 27:72]
  wire  _T_5196 = _T_5195 | _T_5069; // @[Mux.scala 27:72]
  wire  _T_4942 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire  _T_5070 = _T_4942 & way_status_out_42; // @[Mux.scala 27:72]
  wire  _T_5197 = _T_5196 | _T_5070; // @[Mux.scala 27:72]
  wire  _T_4943 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire  _T_5071 = _T_4943 & way_status_out_43; // @[Mux.scala 27:72]
  wire  _T_5198 = _T_5197 | _T_5071; // @[Mux.scala 27:72]
  wire  _T_4944 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire  _T_5072 = _T_4944 & way_status_out_44; // @[Mux.scala 27:72]
  wire  _T_5199 = _T_5198 | _T_5072; // @[Mux.scala 27:72]
  wire  _T_4945 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire  _T_5073 = _T_4945 & way_status_out_45; // @[Mux.scala 27:72]
  wire  _T_5200 = _T_5199 | _T_5073; // @[Mux.scala 27:72]
  wire  _T_4946 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire  _T_5074 = _T_4946 & way_status_out_46; // @[Mux.scala 27:72]
  wire  _T_5201 = _T_5200 | _T_5074; // @[Mux.scala 27:72]
  wire  _T_4947 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire  _T_5075 = _T_4947 & way_status_out_47; // @[Mux.scala 27:72]
  wire  _T_5202 = _T_5201 | _T_5075; // @[Mux.scala 27:72]
  wire  _T_4948 = ifu_ic_rw_int_addr_ff == 7'h30; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire  _T_5076 = _T_4948 & way_status_out_48; // @[Mux.scala 27:72]
  wire  _T_5203 = _T_5202 | _T_5076; // @[Mux.scala 27:72]
  wire  _T_4949 = ifu_ic_rw_int_addr_ff == 7'h31; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire  _T_5077 = _T_4949 & way_status_out_49; // @[Mux.scala 27:72]
  wire  _T_5204 = _T_5203 | _T_5077; // @[Mux.scala 27:72]
  wire  _T_4950 = ifu_ic_rw_int_addr_ff == 7'h32; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire  _T_5078 = _T_4950 & way_status_out_50; // @[Mux.scala 27:72]
  wire  _T_5205 = _T_5204 | _T_5078; // @[Mux.scala 27:72]
  wire  _T_4951 = ifu_ic_rw_int_addr_ff == 7'h33; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire  _T_5079 = _T_4951 & way_status_out_51; // @[Mux.scala 27:72]
  wire  _T_5206 = _T_5205 | _T_5079; // @[Mux.scala 27:72]
  wire  _T_4952 = ifu_ic_rw_int_addr_ff == 7'h34; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire  _T_5080 = _T_4952 & way_status_out_52; // @[Mux.scala 27:72]
  wire  _T_5207 = _T_5206 | _T_5080; // @[Mux.scala 27:72]
  wire  _T_4953 = ifu_ic_rw_int_addr_ff == 7'h35; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire  _T_5081 = _T_4953 & way_status_out_53; // @[Mux.scala 27:72]
  wire  _T_5208 = _T_5207 | _T_5081; // @[Mux.scala 27:72]
  wire  _T_4954 = ifu_ic_rw_int_addr_ff == 7'h36; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire  _T_5082 = _T_4954 & way_status_out_54; // @[Mux.scala 27:72]
  wire  _T_5209 = _T_5208 | _T_5082; // @[Mux.scala 27:72]
  wire  _T_4955 = ifu_ic_rw_int_addr_ff == 7'h37; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire  _T_5083 = _T_4955 & way_status_out_55; // @[Mux.scala 27:72]
  wire  _T_5210 = _T_5209 | _T_5083; // @[Mux.scala 27:72]
  wire  _T_4956 = ifu_ic_rw_int_addr_ff == 7'h38; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire  _T_5084 = _T_4956 & way_status_out_56; // @[Mux.scala 27:72]
  wire  _T_5211 = _T_5210 | _T_5084; // @[Mux.scala 27:72]
  wire  _T_4957 = ifu_ic_rw_int_addr_ff == 7'h39; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire  _T_5085 = _T_4957 & way_status_out_57; // @[Mux.scala 27:72]
  wire  _T_5212 = _T_5211 | _T_5085; // @[Mux.scala 27:72]
  wire  _T_4958 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire  _T_5086 = _T_4958 & way_status_out_58; // @[Mux.scala 27:72]
  wire  _T_5213 = _T_5212 | _T_5086; // @[Mux.scala 27:72]
  wire  _T_4959 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire  _T_5087 = _T_4959 & way_status_out_59; // @[Mux.scala 27:72]
  wire  _T_5214 = _T_5213 | _T_5087; // @[Mux.scala 27:72]
  wire  _T_4960 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire  _T_5088 = _T_4960 & way_status_out_60; // @[Mux.scala 27:72]
  wire  _T_5215 = _T_5214 | _T_5088; // @[Mux.scala 27:72]
  wire  _T_4961 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire  _T_5089 = _T_4961 & way_status_out_61; // @[Mux.scala 27:72]
  wire  _T_5216 = _T_5215 | _T_5089; // @[Mux.scala 27:72]
  wire  _T_4962 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire  _T_5090 = _T_4962 & way_status_out_62; // @[Mux.scala 27:72]
  wire  _T_5217 = _T_5216 | _T_5090; // @[Mux.scala 27:72]
  wire  _T_4963 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire  _T_5091 = _T_4963 & way_status_out_63; // @[Mux.scala 27:72]
  wire  _T_5218 = _T_5217 | _T_5091; // @[Mux.scala 27:72]
  wire  _T_4964 = ifu_ic_rw_int_addr_ff == 7'h40; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire  _T_5092 = _T_4964 & way_status_out_64; // @[Mux.scala 27:72]
  wire  _T_5219 = _T_5218 | _T_5092; // @[Mux.scala 27:72]
  wire  _T_4965 = ifu_ic_rw_int_addr_ff == 7'h41; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire  _T_5093 = _T_4965 & way_status_out_65; // @[Mux.scala 27:72]
  wire  _T_5220 = _T_5219 | _T_5093; // @[Mux.scala 27:72]
  wire  _T_4966 = ifu_ic_rw_int_addr_ff == 7'h42; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire  _T_5094 = _T_4966 & way_status_out_66; // @[Mux.scala 27:72]
  wire  _T_5221 = _T_5220 | _T_5094; // @[Mux.scala 27:72]
  wire  _T_4967 = ifu_ic_rw_int_addr_ff == 7'h43; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire  _T_5095 = _T_4967 & way_status_out_67; // @[Mux.scala 27:72]
  wire  _T_5222 = _T_5221 | _T_5095; // @[Mux.scala 27:72]
  wire  _T_4968 = ifu_ic_rw_int_addr_ff == 7'h44; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire  _T_5096 = _T_4968 & way_status_out_68; // @[Mux.scala 27:72]
  wire  _T_5223 = _T_5222 | _T_5096; // @[Mux.scala 27:72]
  wire  _T_4969 = ifu_ic_rw_int_addr_ff == 7'h45; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire  _T_5097 = _T_4969 & way_status_out_69; // @[Mux.scala 27:72]
  wire  _T_5224 = _T_5223 | _T_5097; // @[Mux.scala 27:72]
  wire  _T_4970 = ifu_ic_rw_int_addr_ff == 7'h46; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire  _T_5098 = _T_4970 & way_status_out_70; // @[Mux.scala 27:72]
  wire  _T_5225 = _T_5224 | _T_5098; // @[Mux.scala 27:72]
  wire  _T_4971 = ifu_ic_rw_int_addr_ff == 7'h47; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire  _T_5099 = _T_4971 & way_status_out_71; // @[Mux.scala 27:72]
  wire  _T_5226 = _T_5225 | _T_5099; // @[Mux.scala 27:72]
  wire  _T_4972 = ifu_ic_rw_int_addr_ff == 7'h48; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire  _T_5100 = _T_4972 & way_status_out_72; // @[Mux.scala 27:72]
  wire  _T_5227 = _T_5226 | _T_5100; // @[Mux.scala 27:72]
  wire  _T_4973 = ifu_ic_rw_int_addr_ff == 7'h49; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire  _T_5101 = _T_4973 & way_status_out_73; // @[Mux.scala 27:72]
  wire  _T_5228 = _T_5227 | _T_5101; // @[Mux.scala 27:72]
  wire  _T_4974 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire  _T_5102 = _T_4974 & way_status_out_74; // @[Mux.scala 27:72]
  wire  _T_5229 = _T_5228 | _T_5102; // @[Mux.scala 27:72]
  wire  _T_4975 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire  _T_5103 = _T_4975 & way_status_out_75; // @[Mux.scala 27:72]
  wire  _T_5230 = _T_5229 | _T_5103; // @[Mux.scala 27:72]
  wire  _T_4976 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire  _T_5104 = _T_4976 & way_status_out_76; // @[Mux.scala 27:72]
  wire  _T_5231 = _T_5230 | _T_5104; // @[Mux.scala 27:72]
  wire  _T_4977 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire  _T_5105 = _T_4977 & way_status_out_77; // @[Mux.scala 27:72]
  wire  _T_5232 = _T_5231 | _T_5105; // @[Mux.scala 27:72]
  wire  _T_4978 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire  _T_5106 = _T_4978 & way_status_out_78; // @[Mux.scala 27:72]
  wire  _T_5233 = _T_5232 | _T_5106; // @[Mux.scala 27:72]
  wire  _T_4979 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire  _T_5107 = _T_4979 & way_status_out_79; // @[Mux.scala 27:72]
  wire  _T_5234 = _T_5233 | _T_5107; // @[Mux.scala 27:72]
  wire  _T_4980 = ifu_ic_rw_int_addr_ff == 7'h50; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire  _T_5108 = _T_4980 & way_status_out_80; // @[Mux.scala 27:72]
  wire  _T_5235 = _T_5234 | _T_5108; // @[Mux.scala 27:72]
  wire  _T_4981 = ifu_ic_rw_int_addr_ff == 7'h51; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire  _T_5109 = _T_4981 & way_status_out_81; // @[Mux.scala 27:72]
  wire  _T_5236 = _T_5235 | _T_5109; // @[Mux.scala 27:72]
  wire  _T_4982 = ifu_ic_rw_int_addr_ff == 7'h52; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire  _T_5110 = _T_4982 & way_status_out_82; // @[Mux.scala 27:72]
  wire  _T_5237 = _T_5236 | _T_5110; // @[Mux.scala 27:72]
  wire  _T_4983 = ifu_ic_rw_int_addr_ff == 7'h53; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire  _T_5111 = _T_4983 & way_status_out_83; // @[Mux.scala 27:72]
  wire  _T_5238 = _T_5237 | _T_5111; // @[Mux.scala 27:72]
  wire  _T_4984 = ifu_ic_rw_int_addr_ff == 7'h54; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire  _T_5112 = _T_4984 & way_status_out_84; // @[Mux.scala 27:72]
  wire  _T_5239 = _T_5238 | _T_5112; // @[Mux.scala 27:72]
  wire  _T_4985 = ifu_ic_rw_int_addr_ff == 7'h55; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire  _T_5113 = _T_4985 & way_status_out_85; // @[Mux.scala 27:72]
  wire  _T_5240 = _T_5239 | _T_5113; // @[Mux.scala 27:72]
  wire  _T_4986 = ifu_ic_rw_int_addr_ff == 7'h56; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire  _T_5114 = _T_4986 & way_status_out_86; // @[Mux.scala 27:72]
  wire  _T_5241 = _T_5240 | _T_5114; // @[Mux.scala 27:72]
  wire  _T_4987 = ifu_ic_rw_int_addr_ff == 7'h57; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire  _T_5115 = _T_4987 & way_status_out_87; // @[Mux.scala 27:72]
  wire  _T_5242 = _T_5241 | _T_5115; // @[Mux.scala 27:72]
  wire  _T_4988 = ifu_ic_rw_int_addr_ff == 7'h58; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire  _T_5116 = _T_4988 & way_status_out_88; // @[Mux.scala 27:72]
  wire  _T_5243 = _T_5242 | _T_5116; // @[Mux.scala 27:72]
  wire  _T_4989 = ifu_ic_rw_int_addr_ff == 7'h59; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire  _T_5117 = _T_4989 & way_status_out_89; // @[Mux.scala 27:72]
  wire  _T_5244 = _T_5243 | _T_5117; // @[Mux.scala 27:72]
  wire  _T_4990 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire  _T_5118 = _T_4990 & way_status_out_90; // @[Mux.scala 27:72]
  wire  _T_5245 = _T_5244 | _T_5118; // @[Mux.scala 27:72]
  wire  _T_4991 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire  _T_5119 = _T_4991 & way_status_out_91; // @[Mux.scala 27:72]
  wire  _T_5246 = _T_5245 | _T_5119; // @[Mux.scala 27:72]
  wire  _T_4992 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire  _T_5120 = _T_4992 & way_status_out_92; // @[Mux.scala 27:72]
  wire  _T_5247 = _T_5246 | _T_5120; // @[Mux.scala 27:72]
  wire  _T_4993 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire  _T_5121 = _T_4993 & way_status_out_93; // @[Mux.scala 27:72]
  wire  _T_5248 = _T_5247 | _T_5121; // @[Mux.scala 27:72]
  wire  _T_4994 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire  _T_5122 = _T_4994 & way_status_out_94; // @[Mux.scala 27:72]
  wire  _T_5249 = _T_5248 | _T_5122; // @[Mux.scala 27:72]
  wire  _T_4995 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire  _T_5123 = _T_4995 & way_status_out_95; // @[Mux.scala 27:72]
  wire  _T_5250 = _T_5249 | _T_5123; // @[Mux.scala 27:72]
  wire  _T_4996 = ifu_ic_rw_int_addr_ff == 7'h60; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire  _T_5124 = _T_4996 & way_status_out_96; // @[Mux.scala 27:72]
  wire  _T_5251 = _T_5250 | _T_5124; // @[Mux.scala 27:72]
  wire  _T_4997 = ifu_ic_rw_int_addr_ff == 7'h61; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire  _T_5125 = _T_4997 & way_status_out_97; // @[Mux.scala 27:72]
  wire  _T_5252 = _T_5251 | _T_5125; // @[Mux.scala 27:72]
  wire  _T_4998 = ifu_ic_rw_int_addr_ff == 7'h62; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire  _T_5126 = _T_4998 & way_status_out_98; // @[Mux.scala 27:72]
  wire  _T_5253 = _T_5252 | _T_5126; // @[Mux.scala 27:72]
  wire  _T_4999 = ifu_ic_rw_int_addr_ff == 7'h63; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire  _T_5127 = _T_4999 & way_status_out_99; // @[Mux.scala 27:72]
  wire  _T_5254 = _T_5253 | _T_5127; // @[Mux.scala 27:72]
  wire  _T_5000 = ifu_ic_rw_int_addr_ff == 7'h64; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire  _T_5128 = _T_5000 & way_status_out_100; // @[Mux.scala 27:72]
  wire  _T_5255 = _T_5254 | _T_5128; // @[Mux.scala 27:72]
  wire  _T_5001 = ifu_ic_rw_int_addr_ff == 7'h65; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire  _T_5129 = _T_5001 & way_status_out_101; // @[Mux.scala 27:72]
  wire  _T_5256 = _T_5255 | _T_5129; // @[Mux.scala 27:72]
  wire  _T_5002 = ifu_ic_rw_int_addr_ff == 7'h66; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire  _T_5130 = _T_5002 & way_status_out_102; // @[Mux.scala 27:72]
  wire  _T_5257 = _T_5256 | _T_5130; // @[Mux.scala 27:72]
  wire  _T_5003 = ifu_ic_rw_int_addr_ff == 7'h67; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire  _T_5131 = _T_5003 & way_status_out_103; // @[Mux.scala 27:72]
  wire  _T_5258 = _T_5257 | _T_5131; // @[Mux.scala 27:72]
  wire  _T_5004 = ifu_ic_rw_int_addr_ff == 7'h68; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire  _T_5132 = _T_5004 & way_status_out_104; // @[Mux.scala 27:72]
  wire  _T_5259 = _T_5258 | _T_5132; // @[Mux.scala 27:72]
  wire  _T_5005 = ifu_ic_rw_int_addr_ff == 7'h69; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire  _T_5133 = _T_5005 & way_status_out_105; // @[Mux.scala 27:72]
  wire  _T_5260 = _T_5259 | _T_5133; // @[Mux.scala 27:72]
  wire  _T_5006 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire  _T_5134 = _T_5006 & way_status_out_106; // @[Mux.scala 27:72]
  wire  _T_5261 = _T_5260 | _T_5134; // @[Mux.scala 27:72]
  wire  _T_5007 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire  _T_5135 = _T_5007 & way_status_out_107; // @[Mux.scala 27:72]
  wire  _T_5262 = _T_5261 | _T_5135; // @[Mux.scala 27:72]
  wire  _T_5008 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire  _T_5136 = _T_5008 & way_status_out_108; // @[Mux.scala 27:72]
  wire  _T_5263 = _T_5262 | _T_5136; // @[Mux.scala 27:72]
  wire  _T_5009 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire  _T_5137 = _T_5009 & way_status_out_109; // @[Mux.scala 27:72]
  wire  _T_5264 = _T_5263 | _T_5137; // @[Mux.scala 27:72]
  wire  _T_5010 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire  _T_5138 = _T_5010 & way_status_out_110; // @[Mux.scala 27:72]
  wire  _T_5265 = _T_5264 | _T_5138; // @[Mux.scala 27:72]
  wire  _T_5011 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire  _T_5139 = _T_5011 & way_status_out_111; // @[Mux.scala 27:72]
  wire  _T_5266 = _T_5265 | _T_5139; // @[Mux.scala 27:72]
  wire  _T_5012 = ifu_ic_rw_int_addr_ff == 7'h70; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire  _T_5140 = _T_5012 & way_status_out_112; // @[Mux.scala 27:72]
  wire  _T_5267 = _T_5266 | _T_5140; // @[Mux.scala 27:72]
  wire  _T_5013 = ifu_ic_rw_int_addr_ff == 7'h71; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire  _T_5141 = _T_5013 & way_status_out_113; // @[Mux.scala 27:72]
  wire  _T_5268 = _T_5267 | _T_5141; // @[Mux.scala 27:72]
  wire  _T_5014 = ifu_ic_rw_int_addr_ff == 7'h72; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire  _T_5142 = _T_5014 & way_status_out_114; // @[Mux.scala 27:72]
  wire  _T_5269 = _T_5268 | _T_5142; // @[Mux.scala 27:72]
  wire  _T_5015 = ifu_ic_rw_int_addr_ff == 7'h73; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire  _T_5143 = _T_5015 & way_status_out_115; // @[Mux.scala 27:72]
  wire  _T_5270 = _T_5269 | _T_5143; // @[Mux.scala 27:72]
  wire  _T_5016 = ifu_ic_rw_int_addr_ff == 7'h74; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire  _T_5144 = _T_5016 & way_status_out_116; // @[Mux.scala 27:72]
  wire  _T_5271 = _T_5270 | _T_5144; // @[Mux.scala 27:72]
  wire  _T_5017 = ifu_ic_rw_int_addr_ff == 7'h75; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire  _T_5145 = _T_5017 & way_status_out_117; // @[Mux.scala 27:72]
  wire  _T_5272 = _T_5271 | _T_5145; // @[Mux.scala 27:72]
  wire  _T_5018 = ifu_ic_rw_int_addr_ff == 7'h76; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire  _T_5146 = _T_5018 & way_status_out_118; // @[Mux.scala 27:72]
  wire  _T_5273 = _T_5272 | _T_5146; // @[Mux.scala 27:72]
  wire  _T_5019 = ifu_ic_rw_int_addr_ff == 7'h77; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire  _T_5147 = _T_5019 & way_status_out_119; // @[Mux.scala 27:72]
  wire  _T_5274 = _T_5273 | _T_5147; // @[Mux.scala 27:72]
  wire  _T_5020 = ifu_ic_rw_int_addr_ff == 7'h78; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire  _T_5148 = _T_5020 & way_status_out_120; // @[Mux.scala 27:72]
  wire  _T_5275 = _T_5274 | _T_5148; // @[Mux.scala 27:72]
  wire  _T_5021 = ifu_ic_rw_int_addr_ff == 7'h79; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire  _T_5149 = _T_5021 & way_status_out_121; // @[Mux.scala 27:72]
  wire  _T_5276 = _T_5275 | _T_5149; // @[Mux.scala 27:72]
  wire  _T_5022 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire  _T_5150 = _T_5022 & way_status_out_122; // @[Mux.scala 27:72]
  wire  _T_5277 = _T_5276 | _T_5150; // @[Mux.scala 27:72]
  wire  _T_5023 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire  _T_5151 = _T_5023 & way_status_out_123; // @[Mux.scala 27:72]
  wire  _T_5278 = _T_5277 | _T_5151; // @[Mux.scala 27:72]
  wire  _T_5024 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire  _T_5152 = _T_5024 & way_status_out_124; // @[Mux.scala 27:72]
  wire  _T_5279 = _T_5278 | _T_5152; // @[Mux.scala 27:72]
  wire  _T_5025 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire  _T_5153 = _T_5025 & way_status_out_125; // @[Mux.scala 27:72]
  wire  _T_5280 = _T_5279 | _T_5153; // @[Mux.scala 27:72]
  wire  _T_5026 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire  _T_5154 = _T_5026 & way_status_out_126; // @[Mux.scala 27:72]
  wire  _T_5281 = _T_5280 | _T_5154; // @[Mux.scala 27:72]
  wire  _T_5027 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[ifu_mem_ctl.scala 628:80]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire  _T_5155 = _T_5027 & way_status_out_127; // @[Mux.scala 27:72]
  wire  way_status = _T_5281 | _T_5155; // @[Mux.scala 27:72]
  wire  _T_198 = ~reset_all_tags; // @[ifu_mem_ctl.scala 164:96]
  wire  _T_200 = _T_198 & _T_339; // @[ifu_mem_ctl.scala 164:112]
  wire [1:0] _T_202 = _T_200 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_203 = _T_202 & io_ic_tag_valid; // @[ifu_mem_ctl.scala 164:135]
  reg [1:0] tagv_mb_scnd_ff; // @[Reg.scala 27:20]
  reg  uncacheable_miss_scnd_ff; // @[Reg.scala 27:20]
  reg [30:0] imb_scnd_ff; // @[Reg.scala 27:20]
  wire [2:0] _T_212 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_212; // @[ifu_mem_ctl.scala 173:45]
  wire  _T_218 = _T_237 | _T_245; // @[ifu_mem_ctl.scala 178:59]
  wire  _T_220 = _T_218 | _T_2274; // @[ifu_mem_ctl.scala 178:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_220; // @[ifu_mem_ctl.scala 178:41]
  wire  _T_225 = _T_233 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 184:39]
  wire  _T_227 = _T_225 & _T_198; // @[ifu_mem_ctl.scala 184:60]
  wire  _T_231 = _T_227 & _T_218; // @[ifu_mem_ctl.scala 184:78]
  wire  ic_act_hit_f = _T_231 & _T_253; // @[ifu_mem_ctl.scala 184:126]
  wire  _T_268 = ic_act_hit_f | ic_byp_hit_f; // @[ifu_mem_ctl.scala 191:31]
  wire  _T_269 = _T_268 | ic_iccm_hit_f; // @[ifu_mem_ctl.scala 191:46]
  wire  _T_270 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 191:94]
  wire  _T_274 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[ifu_mem_ctl.scala 192:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_274; // @[ifu_mem_ctl.scala 192:32]
  wire  _T_280 = imb_ff[11:5] == imb_scnd_ff[11:5]; // @[ifu_mem_ctl.scala 195:79]
  wire  _T_281 = _T_280 & scnd_miss_req; // @[ifu_mem_ctl.scala 195:135]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2737 = |ifu_bus_rresp_ff; // @[ifu_mem_ctl.scala 522:48]
  wire  _T_2738 = _T_2737 & ifu_bus_rvalid_ff; // @[ifu_mem_ctl.scala 522:52]
  wire  bus_ifu_wr_data_error_ff = _T_2738 & miss_pending; // @[ifu_mem_ctl.scala 522:73]
  reg  ifu_wr_data_comb_err_ff; // @[Reg.scala 27:20]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[ifu_mem_ctl.scala 271:59]
  wire  _T_282 = ~ifu_wr_cumulative_err_data; // @[ifu_mem_ctl.scala 195:153]
  wire  scnd_miss_index_match = _T_281 & _T_282; // @[ifu_mem_ctl.scala 195:151]
  wire  _T_283 = ~scnd_miss_index_match; // @[ifu_mem_ctl.scala 198:47]
  wire  _T_284 = scnd_miss_req & _T_283; // @[ifu_mem_ctl.scala 198:45]
  wire  _T_286 = scnd_miss_req & scnd_miss_index_match; // @[ifu_mem_ctl.scala 199:24]
  reg  way_status_mb_ff; // @[Reg.scala 27:20]
  wire  _T_10506 = ~way_status_mb_ff; // @[ifu_mem_ctl.scala 680:31]
  reg [1:0] tagv_mb_ff; // @[Reg.scala 27:20]
  wire  _T_10508 = _T_10506 & tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 680:49]
  wire  _T_10510 = _T_10508 & tagv_mb_ff[1]; // @[ifu_mem_ctl.scala 680:65]
  wire  _T_10512 = ~tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 680:84]
  wire  replace_way_mb_any_0 = _T_10510 | _T_10512; // @[ifu_mem_ctl.scala 680:82]
  wire [1:0] _T_293 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10515 = way_status_mb_ff & tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 681:48]
  wire  _T_10517 = _T_10515 & tagv_mb_ff[1]; // @[ifu_mem_ctl.scala 681:64]
  wire  _T_10519 = ~tagv_mb_ff[1]; // @[ifu_mem_ctl.scala 681:83]
  wire  _T_10521 = _T_10519 & tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 681:98]
  wire  replace_way_mb_any_1 = _T_10517 | _T_10521; // @[ifu_mem_ctl.scala 681:81]
  wire [1:0] _T_294 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_295 = _T_293 & _T_294; // @[ifu_mem_ctl.scala 203:110]
  wire [1:0] _T_296 = tagv_mb_scnd_ff | _T_295; // @[ifu_mem_ctl.scala 203:62]
  wire [1:0] _T_303 = io_ic_tag_valid & _T_202; // @[ifu_mem_ctl.scala 204:58]
  wire  _T_305 = ~scnd_miss_req_q; // @[ifu_mem_ctl.scala 207:36]
  wire  _T_306 = miss_pending & _T_305; // @[ifu_mem_ctl.scala 207:34]
  reg  reset_ic_ff; // @[Reg.scala 27:20]
  wire  _T_307 = reset_all_tags | reset_ic_ff; // @[ifu_mem_ctl.scala 207:72]
  wire  reset_ic_in = _T_306 & _T_307; // @[ifu_mem_ctl.scala 207:53]
  wire  _T_309 = reset_ic_in ^ reset_ic_ff; // @[lib.scala 453:21]
  wire  _T_310 = |_T_309; // @[lib.scala 453:29]
  reg  fetch_uncacheable_ff; // @[Reg.scala 27:20]
  wire  _T_312 = io_ifc_fetch_uncacheable_bf ^ fetch_uncacheable_ff; // @[lib.scala 475:21]
  wire  _T_313 = |_T_312; // @[lib.scala 475:29]
  reg [25:0] miss_addr; // @[Reg.scala 27:20]
  wire  _T_325 = io_ifu_bus_clk_en | ic_act_miss_f; // @[ifu_mem_ctl.scala 219:89]
  wire  _T_326 = _T_325 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 219:105]
  wire  _T_332 = _T_2289 & flush_final_f; // @[ifu_mem_ctl.scala 223:87]
  wire  _T_333 = ~_T_332; // @[ifu_mem_ctl.scala 223:55]
  wire  _T_334 = io_ifc_fetch_req_bf & _T_333; // @[ifu_mem_ctl.scala 223:53]
  wire  _T_2281 = ~_T_2276; // @[ifu_mem_ctl.scala 362:46]
  wire  _T_2282 = _T_2274 & _T_2281; // @[ifu_mem_ctl.scala 362:44]
  wire  stream_miss_f = _T_2282 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 362:84]
  wire  _T_335 = ~stream_miss_f; // @[ifu_mem_ctl.scala 223:106]
  wire  ifc_fetch_req_qual_bf = _T_334 & _T_335; // @[ifu_mem_ctl.scala 223:104]
  wire  _T_336 = ifc_fetch_req_qual_bf ^ ifc_fetch_req_f_raw; // @[lib.scala 475:21]
  wire  _T_337 = |_T_336; // @[lib.scala 475:29]
  wire  _T_10655 = ~io_ifc_iccm_access_bf; // @[ifu_mem_ctl.scala 737:40]
  wire [31:0] _T_10608 = {io_ifc_fetch_addr_bf,1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_10609 = _T_10608 | 32'h7fffffff; // @[ifu_mem_ctl.scala 728:63]
  wire  _T_10611 = _T_10609 == 32'h7fffffff; // @[ifu_mem_ctl.scala 728:94]
  wire [31:0] _T_10615 = _T_10608 | 32'h3fffffff; // @[ifu_mem_ctl.scala 729:63]
  wire  _T_10617 = _T_10615 == 32'hffffffff; // @[ifu_mem_ctl.scala 729:94]
  wire  _T_10619 = _T_10611 | _T_10617; // @[ifu_mem_ctl.scala 728:160]
  wire [31:0] _T_10621 = _T_10608 | 32'h1fffffff; // @[ifu_mem_ctl.scala 730:63]
  wire  _T_10623 = _T_10621 == 32'hbfffffff; // @[ifu_mem_ctl.scala 730:94]
  wire  _T_10625 = _T_10619 | _T_10623; // @[ifu_mem_ctl.scala 729:160]
  wire [31:0] _T_10627 = _T_10608 | 32'hfffffff; // @[ifu_mem_ctl.scala 731:63]
  wire  _T_10629 = _T_10627 == 32'h8fffffff; // @[ifu_mem_ctl.scala 731:94]
  wire  _T_10631 = _T_10625 | _T_10629; // @[ifu_mem_ctl.scala 730:160]
  wire  _T_10637 = _T_10631; // @[ifu_mem_ctl.scala 731:160]
  wire  ifc_region_acc_okay = _T_10631; // @[ifu_mem_ctl.scala 734:160]
  wire  _T_10656 = ~_T_10637; // @[ifu_mem_ctl.scala 737:65]
  wire  _T_10657 = _T_10655 & _T_10656; // @[ifu_mem_ctl.scala 737:63]
  wire  ifc_region_acc_fault_memory_bf = _T_10657 & io_ifc_fetch_req_bf; // @[ifu_mem_ctl.scala 737:86]
  wire  ifc_region_acc_fault_final_bf = io_ifc_region_acc_fault_bf | ifc_region_acc_fault_memory_bf; // @[ifu_mem_ctl.scala 738:63]
  reg  ifc_region_acc_fault_f; // @[Reg.scala 27:20]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_345 = _T_245 | _T_2274; // @[ifu_mem_ctl.scala 231:55]
  wire  _T_348 = _T_345 & _T_59; // @[ifu_mem_ctl.scala 231:82]
  wire  _T_2295 = ~ifu_bus_rid_ff[0]; // @[ifu_mem_ctl.scala 367:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2295}; // @[Cat.scala 29:58]
  wire  _T_2296 = other_tag == 3'h0; // @[ifu_mem_ctl.scala 368:81]
  wire  _T_2320 = _T_2296 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2299 = other_tag == 3'h1; // @[ifu_mem_ctl.scala 368:81]
  wire  _T_2321 = _T_2299 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2328 = _T_2320 | _T_2321; // @[Mux.scala 27:72]
  wire  _T_2302 = other_tag == 3'h2; // @[ifu_mem_ctl.scala 368:81]
  wire  _T_2322 = _T_2302 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2329 = _T_2328 | _T_2322; // @[Mux.scala 27:72]
  wire  _T_2305 = other_tag == 3'h3; // @[ifu_mem_ctl.scala 368:81]
  wire  _T_2323 = _T_2305 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2330 = _T_2329 | _T_2323; // @[Mux.scala 27:72]
  wire  _T_2308 = other_tag == 3'h4; // @[ifu_mem_ctl.scala 368:81]
  wire  _T_2324 = _T_2308 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2331 = _T_2330 | _T_2324; // @[Mux.scala 27:72]
  wire  _T_2311 = other_tag == 3'h5; // @[ifu_mem_ctl.scala 368:81]
  wire  _T_2325 = _T_2311 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2332 = _T_2331 | _T_2325; // @[Mux.scala 27:72]
  wire  _T_2314 = other_tag == 3'h6; // @[ifu_mem_ctl.scala 368:81]
  wire  _T_2326 = _T_2314 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2333 = _T_2332 | _T_2326; // @[Mux.scala 27:72]
  wire  _T_2317 = other_tag == 3'h7; // @[ifu_mem_ctl.scala 368:81]
  wire  _T_2327 = _T_2317 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2333 | _T_2327; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[ifu_mem_ctl.scala 369:46]
  wire  _T_352 = miss_pending & write_ic_16_bytes; // @[ifu_mem_ctl.scala 235:35]
  wire  _T_354 = _T_352 & _T_20; // @[ifu_mem_ctl.scala 235:55]
  reg  ic_act_miss_f_delayed; // @[Reg.scala 27:20]
  wire  _T_2731 = ic_act_miss_f_delayed & _T_2290; // @[ifu_mem_ctl.scala 520:53]
  wire  reset_tag_valid_for_miss = _T_2731 & _T_20; // @[ifu_mem_ctl.scala 520:84]
  wire  sel_mb_addr = _T_354 | reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 235:79]
  wire [30:0] _T_358 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_359 = ~sel_mb_addr; // @[ifu_mem_ctl.scala 237:5]
  wire [30:0] _T_360 = sel_mb_addr ? _T_358 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_361 = _T_359 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire  _T_367 = _T_354 & last_beat; // @[ifu_mem_ctl.scala 239:85]
  wire  _T_2722 = ~_T_2737; // @[ifu_mem_ctl.scala 517:84]
  wire  _T_2723 = _T_103 & _T_2722; // @[ifu_mem_ctl.scala 517:82]
  wire  bus_ifu_wr_en_ff_q = _T_2723 & write_ic_16_bytes; // @[ifu_mem_ctl.scala 517:108]
  wire  _T_368 = _T_367 & bus_ifu_wr_en_ff_q; // @[ifu_mem_ctl.scala 239:97]
  wire  sel_mb_status_addr = _T_368 | reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 239:119]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_358 : ifu_fetch_addr_int_f; // @[ifu_mem_ctl.scala 240:31]
  wire  _T_374 = sel_mb_addr ^ sel_mb_addr_ff; // @[lib.scala 475:21]
  wire  _T_375 = |_T_374; // @[lib.scala 475:29]
  wire  _T_377 = io_ifu_bus_clk_en & io_ifu_axi_r_valid; // @[ifu_mem_ctl.scala 242:74]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] _T_595 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[lib.scala 276:13]
  wire  _T_596 = ^_T_595; // @[lib.scala 276:20]
  wire [6:0] _T_602 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[lib.scala 276:30]
  wire [7:0] _T_609 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[lib.scala 276:30]
  wire [14:0] _T_610 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_602}; // @[lib.scala 276:30]
  wire [7:0] _T_617 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[lib.scala 276:30]
  wire [30:0] _T_626 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_617,_T_610}; // @[lib.scala 276:30]
  wire  _T_627 = ^_T_626; // @[lib.scala 276:37]
  wire [6:0] _T_633 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[lib.scala 276:47]
  wire [14:0] _T_641 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_633}; // @[lib.scala 276:47]
  wire [30:0] _T_657 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_617,_T_641}; // @[lib.scala 276:47]
  wire  _T_658 = ^_T_657; // @[lib.scala 276:54]
  wire [6:0] _T_664 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[lib.scala 276:64]
  wire [14:0] _T_672 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_664}; // @[lib.scala 276:64]
  wire [30:0] _T_688 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_609,_T_672}; // @[lib.scala 276:64]
  wire  _T_689 = ^_T_688; // @[lib.scala 276:71]
  wire [7:0] _T_696 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[lib.scala 276:81]
  wire [16:0] _T_705 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_696}; // @[lib.scala 276:81]
  wire [8:0] _T_713 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[lib.scala 276:81]
  wire [17:0] _T_722 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_713}; // @[lib.scala 276:81]
  wire [34:0] _T_723 = {_T_722,_T_705}; // @[lib.scala 276:81]
  wire  _T_724 = ^_T_723; // @[lib.scala 276:88]
  wire [7:0] _T_731 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[lib.scala 276:98]
  wire [16:0] _T_740 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_731}; // @[lib.scala 276:98]
  wire [8:0] _T_748 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[lib.scala 276:98]
  wire [17:0] _T_757 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_748}; // @[lib.scala 276:98]
  wire [34:0] _T_758 = {_T_757,_T_740}; // @[lib.scala 276:98]
  wire  _T_759 = ^_T_758; // @[lib.scala 276:105]
  wire [7:0] _T_766 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[lib.scala 276:115]
  wire [16:0] _T_775 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_766}; // @[lib.scala 276:115]
  wire [8:0] _T_783 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[lib.scala 276:115]
  wire [17:0] _T_792 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_783}; // @[lib.scala 276:115]
  wire [34:0] _T_793 = {_T_792,_T_775}; // @[lib.scala 276:115]
  wire  _T_794 = ^_T_793; // @[lib.scala 276:122]
  wire [3:0] _T_2336 = {ifu_bus_rid_ff[2:1],_T_2295,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2337 = _T_2336 == 4'h0; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_2384 = _T_2337 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2340 = _T_2336 == 4'h1; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_2385 = _T_2340 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2400 = _T_2384 | _T_2385; // @[Mux.scala 27:72]
  wire  _T_2343 = _T_2336 == 4'h2; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_2386 = _T_2343 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2401 = _T_2400 | _T_2386; // @[Mux.scala 27:72]
  wire  _T_2346 = _T_2336 == 4'h3; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_2387 = _T_2346 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2402 = _T_2401 | _T_2387; // @[Mux.scala 27:72]
  wire  _T_2349 = _T_2336 == 4'h4; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_2388 = _T_2349 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2403 = _T_2402 | _T_2388; // @[Mux.scala 27:72]
  wire  _T_2352 = _T_2336 == 4'h5; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_2389 = _T_2352 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2404 = _T_2403 | _T_2389; // @[Mux.scala 27:72]
  wire  _T_2355 = _T_2336 == 4'h6; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_2390 = _T_2355 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2405 = _T_2404 | _T_2390; // @[Mux.scala 27:72]
  wire  _T_2358 = _T_2336 == 4'h7; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_2391 = _T_2358 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2406 = _T_2405 | _T_2391; // @[Mux.scala 27:72]
  wire  _T_2361 = _T_2336 == 4'h8; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_2392 = _T_2361 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2407 = _T_2406 | _T_2392; // @[Mux.scala 27:72]
  wire  _T_2364 = _T_2336 == 4'h9; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_2393 = _T_2364 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2408 = _T_2407 | _T_2393; // @[Mux.scala 27:72]
  wire  _T_2367 = _T_2336 == 4'ha; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_2394 = _T_2367 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2409 = _T_2408 | _T_2394; // @[Mux.scala 27:72]
  wire  _T_2370 = _T_2336 == 4'hb; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_2395 = _T_2370 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2410 = _T_2409 | _T_2395; // @[Mux.scala 27:72]
  wire  _T_2373 = _T_2336 == 4'hc; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_2396 = _T_2373 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2411 = _T_2410 | _T_2396; // @[Mux.scala 27:72]
  wire  _T_2376 = _T_2336 == 4'hd; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_2397 = _T_2376 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2412 = _T_2411 | _T_2397; // @[Mux.scala 27:72]
  wire  _T_2379 = _T_2336 == 4'he; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_2398 = _T_2379 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2413 = _T_2412 | _T_2398; // @[Mux.scala 27:72]
  wire  _T_2382 = _T_2336 == 4'hf; // @[ifu_mem_ctl.scala 370:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_2399 = _T_2382 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2414 = _T_2413 | _T_2399; // @[Mux.scala 27:72]
  wire [3:0] _T_2416 = {ifu_bus_rid_ff[2:1],_T_2295,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2417 = _T_2416 == 4'h0; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2464 = _T_2417 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2420 = _T_2416 == 4'h1; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2465 = _T_2420 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2480 = _T_2464 | _T_2465; // @[Mux.scala 27:72]
  wire  _T_2423 = _T_2416 == 4'h2; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2466 = _T_2423 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2481 = _T_2480 | _T_2466; // @[Mux.scala 27:72]
  wire  _T_2426 = _T_2416 == 4'h3; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2467 = _T_2426 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2482 = _T_2481 | _T_2467; // @[Mux.scala 27:72]
  wire  _T_2429 = _T_2416 == 4'h4; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2468 = _T_2429 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2483 = _T_2482 | _T_2468; // @[Mux.scala 27:72]
  wire  _T_2432 = _T_2416 == 4'h5; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2469 = _T_2432 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2484 = _T_2483 | _T_2469; // @[Mux.scala 27:72]
  wire  _T_2435 = _T_2416 == 4'h6; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2470 = _T_2435 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2485 = _T_2484 | _T_2470; // @[Mux.scala 27:72]
  wire  _T_2438 = _T_2416 == 4'h7; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2471 = _T_2438 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2486 = _T_2485 | _T_2471; // @[Mux.scala 27:72]
  wire  _T_2441 = _T_2416 == 4'h8; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2472 = _T_2441 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2487 = _T_2486 | _T_2472; // @[Mux.scala 27:72]
  wire  _T_2444 = _T_2416 == 4'h9; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2473 = _T_2444 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2488 = _T_2487 | _T_2473; // @[Mux.scala 27:72]
  wire  _T_2447 = _T_2416 == 4'ha; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2474 = _T_2447 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2489 = _T_2488 | _T_2474; // @[Mux.scala 27:72]
  wire  _T_2450 = _T_2416 == 4'hb; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2475 = _T_2450 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2490 = _T_2489 | _T_2475; // @[Mux.scala 27:72]
  wire  _T_2453 = _T_2416 == 4'hc; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2476 = _T_2453 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2491 = _T_2490 | _T_2476; // @[Mux.scala 27:72]
  wire  _T_2456 = _T_2416 == 4'hd; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2477 = _T_2456 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2492 = _T_2491 | _T_2477; // @[Mux.scala 27:72]
  wire  _T_2459 = _T_2416 == 4'he; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2478 = _T_2459 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2493 = _T_2492 | _T_2478; // @[Mux.scala 27:72]
  wire  _T_2462 = _T_2416 == 4'hf; // @[ifu_mem_ctl.scala 371:66]
  wire [31:0] _T_2479 = _T_2462 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2494 = _T_2493 | _T_2479; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2414,_T_2494}; // @[Cat.scala 29:58]
  wire [6:0] _T_1017 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[lib.scala 276:13]
  wire  _T_1018 = ^_T_1017; // @[lib.scala 276:20]
  wire [6:0] _T_1024 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[lib.scala 276:30]
  wire [7:0] _T_1031 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[lib.scala 276:30]
  wire [14:0] _T_1032 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_1024}; // @[lib.scala 276:30]
  wire [7:0] _T_1039 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[lib.scala 276:30]
  wire [30:0] _T_1048 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1039,_T_1032}; // @[lib.scala 276:30]
  wire  _T_1049 = ^_T_1048; // @[lib.scala 276:37]
  wire [6:0] _T_1055 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[lib.scala 276:47]
  wire [14:0] _T_1063 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1055}; // @[lib.scala 276:47]
  wire [30:0] _T_1079 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1039,_T_1063}; // @[lib.scala 276:47]
  wire  _T_1080 = ^_T_1079; // @[lib.scala 276:54]
  wire [6:0] _T_1086 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[lib.scala 276:64]
  wire [14:0] _T_1094 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1086}; // @[lib.scala 276:64]
  wire [30:0] _T_1110 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1031,_T_1094}; // @[lib.scala 276:64]
  wire  _T_1111 = ^_T_1110; // @[lib.scala 276:71]
  wire [7:0] _T_1118 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[lib.scala 276:81]
  wire [16:0] _T_1127 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1118}; // @[lib.scala 276:81]
  wire [8:0] _T_1135 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[lib.scala 276:81]
  wire [17:0] _T_1144 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1135}; // @[lib.scala 276:81]
  wire [34:0] _T_1145 = {_T_1144,_T_1127}; // @[lib.scala 276:81]
  wire  _T_1146 = ^_T_1145; // @[lib.scala 276:88]
  wire [7:0] _T_1153 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[lib.scala 276:98]
  wire [16:0] _T_1162 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1153}; // @[lib.scala 276:98]
  wire [8:0] _T_1170 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[lib.scala 276:98]
  wire [17:0] _T_1179 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1170}; // @[lib.scala 276:98]
  wire [34:0] _T_1180 = {_T_1179,_T_1162}; // @[lib.scala 276:98]
  wire  _T_1181 = ^_T_1180; // @[lib.scala 276:105]
  wire [7:0] _T_1188 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[lib.scala 276:115]
  wire [16:0] _T_1197 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1188}; // @[lib.scala 276:115]
  wire [8:0] _T_1205 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[lib.scala 276:115]
  wire [17:0] _T_1214 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1205}; // @[lib.scala 276:115]
  wire [34:0] _T_1215 = {_T_1214,_T_1197}; // @[lib.scala 276:115]
  wire  _T_1216 = ^_T_1215; // @[lib.scala 276:122]
  wire [70:0] _T_1261 = {_T_596,_T_627,_T_658,_T_689,_T_724,_T_759,_T_794,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1260 = {_T_1018,_T_1049,_T_1080,_T_1111,_T_1146,_T_1181,_T_1216,_T_2414,_T_2494}; // @[Cat.scala 29:58]
  wire [141:0] _T_1262 = {_T_596,_T_627,_T_658,_T_689,_T_724,_T_759,_T_794,ifu_bus_rdata_ff,_T_1260}; // @[Cat.scala 29:58]
  wire [141:0] _T_1265 = {_T_1018,_T_1049,_T_1080,_T_1111,_T_1146,_T_1181,_T_1216,_T_2414,_T_2494,_T_1261}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1262 : _T_1265; // @[ifu_mem_ctl.scala 264:28]
  wire  _T_1224 = |io_ic_eccerr; // @[ifu_mem_ctl.scala 252:73]
  wire  _T_1225 = _T_1224 & ic_act_hit_f; // @[ifu_mem_ctl.scala 252:100]
  wire  _T_2498 = io_ic_tag_perr & _T_339; // @[ifu_mem_ctl.scala 374:44]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[ifu_mem_ctl.scala 318:28]
  wire  _T_1436 = bypass_index[4:2] == 3'h0; // @[ifu_mem_ctl.scala 320:114]
  wire  bus_ifu_wr_en = _T_16 & miss_pending; // @[ifu_mem_ctl.scala 515:35]
  wire  _T_1321 = io_ifu_axi_r_bits_id == 3'h0; // @[ifu_mem_ctl.scala 301:96]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1321; // @[ifu_mem_ctl.scala 301:73]
  wire  _T_1362 = ~ic_act_miss_f; // @[ifu_mem_ctl.scala 309:118]
  wire  _T_1363 = ic_miss_buff_data_valid[0] & _T_1362; // @[ifu_mem_ctl.scala 309:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1363; // @[ifu_mem_ctl.scala 309:88]
  wire  _T_1459 = _T_1436 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1439 = bypass_index[4:2] == 3'h1; // @[ifu_mem_ctl.scala 320:114]
  wire  _T_1322 = io_ifu_axi_r_bits_id == 3'h1; // @[ifu_mem_ctl.scala 301:96]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1322; // @[ifu_mem_ctl.scala 301:73]
  wire  _T_1366 = ic_miss_buff_data_valid[1] & _T_1362; // @[ifu_mem_ctl.scala 309:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1366; // @[ifu_mem_ctl.scala 309:88]
  wire  _T_1460 = _T_1439 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1467 = _T_1459 | _T_1460; // @[Mux.scala 27:72]
  wire  _T_1442 = bypass_index[4:2] == 3'h2; // @[ifu_mem_ctl.scala 320:114]
  wire  _T_1323 = io_ifu_axi_r_bits_id == 3'h2; // @[ifu_mem_ctl.scala 301:96]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1323; // @[ifu_mem_ctl.scala 301:73]
  wire  _T_1369 = ic_miss_buff_data_valid[2] & _T_1362; // @[ifu_mem_ctl.scala 309:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1369; // @[ifu_mem_ctl.scala 309:88]
  wire  _T_1461 = _T_1442 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1468 = _T_1467 | _T_1461; // @[Mux.scala 27:72]
  wire  _T_1445 = bypass_index[4:2] == 3'h3; // @[ifu_mem_ctl.scala 320:114]
  wire  _T_1324 = io_ifu_axi_r_bits_id == 3'h3; // @[ifu_mem_ctl.scala 301:96]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1324; // @[ifu_mem_ctl.scala 301:73]
  wire  _T_1372 = ic_miss_buff_data_valid[3] & _T_1362; // @[ifu_mem_ctl.scala 309:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1372; // @[ifu_mem_ctl.scala 309:88]
  wire  _T_1462 = _T_1445 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1469 = _T_1468 | _T_1462; // @[Mux.scala 27:72]
  wire  _T_1448 = bypass_index[4:2] == 3'h4; // @[ifu_mem_ctl.scala 320:114]
  wire  _T_1325 = io_ifu_axi_r_bits_id == 3'h4; // @[ifu_mem_ctl.scala 301:96]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1325; // @[ifu_mem_ctl.scala 301:73]
  wire  _T_1375 = ic_miss_buff_data_valid[4] & _T_1362; // @[ifu_mem_ctl.scala 309:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1375; // @[ifu_mem_ctl.scala 309:88]
  wire  _T_1463 = _T_1448 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1470 = _T_1469 | _T_1463; // @[Mux.scala 27:72]
  wire  _T_1451 = bypass_index[4:2] == 3'h5; // @[ifu_mem_ctl.scala 320:114]
  wire  _T_1326 = io_ifu_axi_r_bits_id == 3'h5; // @[ifu_mem_ctl.scala 301:96]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1326; // @[ifu_mem_ctl.scala 301:73]
  wire  _T_1378 = ic_miss_buff_data_valid[5] & _T_1362; // @[ifu_mem_ctl.scala 309:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1378; // @[ifu_mem_ctl.scala 309:88]
  wire  _T_1464 = _T_1451 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1471 = _T_1470 | _T_1464; // @[Mux.scala 27:72]
  wire  _T_1454 = bypass_index[4:2] == 3'h6; // @[ifu_mem_ctl.scala 320:114]
  wire  _T_1327 = io_ifu_axi_r_bits_id == 3'h6; // @[ifu_mem_ctl.scala 301:96]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1327; // @[ifu_mem_ctl.scala 301:73]
  wire  _T_1381 = ic_miss_buff_data_valid[6] & _T_1362; // @[ifu_mem_ctl.scala 309:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1381; // @[ifu_mem_ctl.scala 309:88]
  wire  _T_1465 = _T_1454 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1472 = _T_1471 | _T_1465; // @[Mux.scala 27:72]
  wire  _T_1457 = bypass_index[4:2] == 3'h7; // @[ifu_mem_ctl.scala 320:114]
  wire  _T_1328 = io_ifu_axi_r_bits_id == 3'h7; // @[ifu_mem_ctl.scala 301:96]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1328; // @[ifu_mem_ctl.scala 301:73]
  wire  _T_1384 = ic_miss_buff_data_valid[7] & _T_1362; // @[ifu_mem_ctl.scala 309:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1384; // @[ifu_mem_ctl.scala 309:88]
  wire  _T_1466 = _T_1457 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1472 | _T_1466; // @[Mux.scala 27:72]
  wire  _T_1475 = ~bypass_index[1]; // @[ifu_mem_ctl.scala 321:58]
  wire  _T_1476 = bypass_valid_value_check & _T_1475; // @[ifu_mem_ctl.scala 321:56]
  wire  _T_1478 = ~bypass_index[0]; // @[ifu_mem_ctl.scala 321:77]
  wire  _T_1479 = _T_1476 & _T_1478; // @[ifu_mem_ctl.scala 321:75]
  wire  _T_1484 = _T_1476 & bypass_index[0]; // @[ifu_mem_ctl.scala 322:50]
  wire  _T_1485 = _T_1479 | _T_1484; // @[ifu_mem_ctl.scala 321:95]
  wire  _T_1487 = bypass_valid_value_check & bypass_index[1]; // @[ifu_mem_ctl.scala 323:31]
  wire  _T_1490 = _T_1487 & _T_1478; // @[ifu_mem_ctl.scala 323:49]
  wire  _T_1491 = _T_1485 | _T_1490; // @[ifu_mem_ctl.scala 322:69]
  wire  _T_1495 = _T_1487 & bypass_index[0]; // @[ifu_mem_ctl.scala 324:49]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[ifu_mem_ctl.scala 319:70]
  wire  _T_1496 = bypass_index_5_3_inc == 3'h0; // @[ifu_mem_ctl.scala 324:130]
  wire  _T_1512 = _T_1496 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1498 = bypass_index_5_3_inc == 3'h1; // @[ifu_mem_ctl.scala 324:130]
  wire  _T_1513 = _T_1498 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1520 = _T_1512 | _T_1513; // @[Mux.scala 27:72]
  wire  _T_1500 = bypass_index_5_3_inc == 3'h2; // @[ifu_mem_ctl.scala 324:130]
  wire  _T_1514 = _T_1500 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1521 = _T_1520 | _T_1514; // @[Mux.scala 27:72]
  wire  _T_1502 = bypass_index_5_3_inc == 3'h3; // @[ifu_mem_ctl.scala 324:130]
  wire  _T_1515 = _T_1502 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1522 = _T_1521 | _T_1515; // @[Mux.scala 27:72]
  wire  _T_1504 = bypass_index_5_3_inc == 3'h4; // @[ifu_mem_ctl.scala 324:130]
  wire  _T_1516 = _T_1504 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1523 = _T_1522 | _T_1516; // @[Mux.scala 27:72]
  wire  _T_1506 = bypass_index_5_3_inc == 3'h5; // @[ifu_mem_ctl.scala 324:130]
  wire  _T_1517 = _T_1506 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1524 = _T_1523 | _T_1517; // @[Mux.scala 27:72]
  wire  _T_1508 = bypass_index_5_3_inc == 3'h6; // @[ifu_mem_ctl.scala 324:130]
  wire  _T_1518 = _T_1508 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1525 = _T_1524 | _T_1518; // @[Mux.scala 27:72]
  wire  _T_1510 = bypass_index_5_3_inc == 3'h7; // @[ifu_mem_ctl.scala 324:130]
  wire  _T_1519 = _T_1510 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1526 = _T_1525 | _T_1519; // @[Mux.scala 27:72]
  wire  _T_1528 = _T_1495 & _T_1526; // @[ifu_mem_ctl.scala 324:67]
  wire  _T_1529 = _T_1491 | _T_1528; // @[ifu_mem_ctl.scala 323:69]
  wire [4:0] _GEN_516 = {{2'd0}, bypass_index[4:2]}; // @[ifu_mem_ctl.scala 325:70]
  wire  _T_1532 = _GEN_516 == 5'h1f; // @[ifu_mem_ctl.scala 325:70]
  wire  _T_1533 = bypass_valid_value_check & _T_1532; // @[ifu_mem_ctl.scala 325:31]
  wire  bypass_data_ready_in = _T_1529 | _T_1533; // @[ifu_mem_ctl.scala 324:179]
  wire  _T_1534 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[ifu_mem_ctl.scala 329:53]
  wire  _T_1535 = _T_1534 & uncacheable_miss_ff; // @[ifu_mem_ctl.scala 329:73]
  wire  _T_1537 = _T_1535 & _T_339; // @[ifu_mem_ctl.scala 329:96]
  wire  _T_1539 = _T_1537 & _T_61; // @[ifu_mem_ctl.scala 329:118]
  wire  _T_1541 = crit_wd_byp_ok_ff & _T_20; // @[ifu_mem_ctl.scala 330:47]
  wire  _T_1543 = _T_1541 & _T_339; // @[ifu_mem_ctl.scala 330:70]
  wire  _T_1545 = _T_1543 & _T_61; // @[ifu_mem_ctl.scala 330:92]
  wire  _T_1546 = _T_1539 | _T_1545; // @[ifu_mem_ctl.scala 329:143]
  reg  ic_crit_wd_rdy_new_ff; // @[Reg.scala 27:20]
  wire  _T_1547 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[ifu_mem_ctl.scala 331:28]
  wire  _T_1548 = ~fetch_req_icache_f; // @[ifu_mem_ctl.scala 331:50]
  wire  _T_1549 = _T_1547 & _T_1548; // @[ifu_mem_ctl.scala 331:48]
  wire  _T_1551 = _T_1549 & _T_339; // @[ifu_mem_ctl.scala 331:70]
  wire  ic_crit_wd_rdy_new_in = _T_1546 | _T_1551; // @[ifu_mem_ctl.scala 330:117]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[ifu_mem_ctl.scala 525:43]
  wire  _T_1278 = ic_crit_wd_rdy | _T_2274; // @[ifu_mem_ctl.scala 276:38]
  wire  _T_1280 = _T_1278 | _T_2290; // @[ifu_mem_ctl.scala 276:64]
  wire  _T_1281 = miss_state == 3'h3; // @[ifu_mem_ctl.scala 276:109]
  wire  _T_1282 = _T_1280 | _T_1281; // @[ifu_mem_ctl.scala 276:95]
  wire  _T_1283 = ~_T_1282; // @[ifu_mem_ctl.scala 276:21]
  wire  _T_1284 = ~fetch_req_iccm_f; // @[ifu_mem_ctl.scala 276:129]
  wire  _T_1285 = _T_1283 & _T_1284; // @[ifu_mem_ctl.scala 276:127]
  wire  sel_ic_data = _T_1285 & _T_215; // @[ifu_mem_ctl.scala 276:147]
  wire  _T_2499 = _T_2498 & sel_ic_data; // @[ifu_mem_ctl.scala 374:66]
  wire [1:0] _T_1298 = ic_byp_hit_f ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg [7:0] ic_miss_buff_data_error; // @[ifu_mem_ctl.scala 315:62]
  wire [7:0] _T_1647 = ic_miss_buff_data_error >> byp_fetch_index[4:2]; // @[ifu_mem_ctl.scala 342:55]
  wire  _T_1651 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 343:34]
  wire  _T_1655 = ~_T_1647[0]; // @[ifu_mem_ctl.scala 343:63]
  wire  _T_1656 = _T_1651 & _T_1655; // @[ifu_mem_ctl.scala 343:61]
  wire [7:0] _T_1658 = ic_miss_buff_data_error >> byp_fetch_index_inc; // @[ifu_mem_ctl.scala 344:46]
  wire  _T_1660 = _T_2275 & _T_1658[0]; // @[ifu_mem_ctl.scala 344:21]
  wire  _T_1661 = _T_1656 & _T_1660; // @[ifu_mem_ctl.scala 343:132]
  wire [1:0] _T_1662 = _T_1661 ? 2'h2 : 2'h0; // @[ifu_mem_ctl.scala 343:8]
  wire [1:0] ifu_byp_data_err_f = _T_1647[0] ? 2'h3 : _T_1662; // @[ifu_mem_ctl.scala 342:31]
  wire [1:0] ifc_bus_acc_fault_f = _T_1298 & ifu_byp_data_err_f; // @[ifu_mem_ctl.scala 289:50]
  wire  _T_2500 = |ifc_bus_acc_fault_f; // @[ifu_mem_ctl.scala 374:136]
  wire  _T_2501 = ifc_region_acc_fault_final_f | _T_2500; // @[ifu_mem_ctl.scala 374:113]
  wire  _T_2502 = ~_T_2501; // @[ifu_mem_ctl.scala 374:82]
  wire  _T_2503 = _T_2499 & _T_2502; // @[ifu_mem_ctl.scala 374:80]
  wire  _T_2505 = fetch_req_icache_f & _T_198; // @[ifu_mem_ctl.scala 375:25]
  wire  _T_2509 = _T_2505 & _T_218; // @[ifu_mem_ctl.scala 375:43]
  wire  _T_2511 = _T_2509 & _T_253; // @[ifu_mem_ctl.scala 375:91]
  wire  ic_rd_parity_final_err = _T_2503 & _T_2511; // @[ifu_mem_ctl.scala 374:142]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_10124 = _T_4900 & ic_tag_valid_out_1_0; // @[ifu_mem_ctl.scala 656:8]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_10126 = _T_4901 & ic_tag_valid_out_1_1; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10379 = _T_10124 | _T_10126; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_10128 = _T_4902 & ic_tag_valid_out_1_2; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10380 = _T_10379 | _T_10128; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_10130 = _T_4903 & ic_tag_valid_out_1_3; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10381 = _T_10380 | _T_10130; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_10132 = _T_4904 & ic_tag_valid_out_1_4; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10382 = _T_10381 | _T_10132; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_10134 = _T_4905 & ic_tag_valid_out_1_5; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10383 = _T_10382 | _T_10134; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_10136 = _T_4906 & ic_tag_valid_out_1_6; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10384 = _T_10383 | _T_10136; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_10138 = _T_4907 & ic_tag_valid_out_1_7; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10385 = _T_10384 | _T_10138; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_10140 = _T_4908 & ic_tag_valid_out_1_8; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10386 = _T_10385 | _T_10140; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_10142 = _T_4909 & ic_tag_valid_out_1_9; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10387 = _T_10386 | _T_10142; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_10144 = _T_4910 & ic_tag_valid_out_1_10; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10388 = _T_10387 | _T_10144; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_10146 = _T_4911 & ic_tag_valid_out_1_11; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10389 = _T_10388 | _T_10146; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_10148 = _T_4912 & ic_tag_valid_out_1_12; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10390 = _T_10389 | _T_10148; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_10150 = _T_4913 & ic_tag_valid_out_1_13; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10391 = _T_10390 | _T_10150; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_10152 = _T_4914 & ic_tag_valid_out_1_14; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10392 = _T_10391 | _T_10152; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_10154 = _T_4915 & ic_tag_valid_out_1_15; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10393 = _T_10392 | _T_10154; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_10156 = _T_4916 & ic_tag_valid_out_1_16; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10394 = _T_10393 | _T_10156; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_10158 = _T_4917 & ic_tag_valid_out_1_17; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10395 = _T_10394 | _T_10158; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_10160 = _T_4918 & ic_tag_valid_out_1_18; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10396 = _T_10395 | _T_10160; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_10162 = _T_4919 & ic_tag_valid_out_1_19; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10397 = _T_10396 | _T_10162; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_10164 = _T_4920 & ic_tag_valid_out_1_20; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10398 = _T_10397 | _T_10164; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_10166 = _T_4921 & ic_tag_valid_out_1_21; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10399 = _T_10398 | _T_10166; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_10168 = _T_4922 & ic_tag_valid_out_1_22; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10400 = _T_10399 | _T_10168; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_10170 = _T_4923 & ic_tag_valid_out_1_23; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10401 = _T_10400 | _T_10170; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_10172 = _T_4924 & ic_tag_valid_out_1_24; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10402 = _T_10401 | _T_10172; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_10174 = _T_4925 & ic_tag_valid_out_1_25; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10403 = _T_10402 | _T_10174; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_10176 = _T_4926 & ic_tag_valid_out_1_26; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10404 = _T_10403 | _T_10176; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_10178 = _T_4927 & ic_tag_valid_out_1_27; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10405 = _T_10404 | _T_10178; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_10180 = _T_4928 & ic_tag_valid_out_1_28; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10406 = _T_10405 | _T_10180; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_10182 = _T_4929 & ic_tag_valid_out_1_29; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10407 = _T_10406 | _T_10182; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_10184 = _T_4930 & ic_tag_valid_out_1_30; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10408 = _T_10407 | _T_10184; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_10186 = _T_4931 & ic_tag_valid_out_1_31; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10409 = _T_10408 | _T_10186; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_10188 = _T_4932 & ic_tag_valid_out_1_32; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10410 = _T_10409 | _T_10188; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_10190 = _T_4933 & ic_tag_valid_out_1_33; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10411 = _T_10410 | _T_10190; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_10192 = _T_4934 & ic_tag_valid_out_1_34; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10412 = _T_10411 | _T_10192; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_10194 = _T_4935 & ic_tag_valid_out_1_35; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10413 = _T_10412 | _T_10194; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_10196 = _T_4936 & ic_tag_valid_out_1_36; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10414 = _T_10413 | _T_10196; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_10198 = _T_4937 & ic_tag_valid_out_1_37; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10415 = _T_10414 | _T_10198; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_10200 = _T_4938 & ic_tag_valid_out_1_38; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10416 = _T_10415 | _T_10200; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_10202 = _T_4939 & ic_tag_valid_out_1_39; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10417 = _T_10416 | _T_10202; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_10204 = _T_4940 & ic_tag_valid_out_1_40; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10418 = _T_10417 | _T_10204; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_10206 = _T_4941 & ic_tag_valid_out_1_41; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10419 = _T_10418 | _T_10206; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_10208 = _T_4942 & ic_tag_valid_out_1_42; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10420 = _T_10419 | _T_10208; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_10210 = _T_4943 & ic_tag_valid_out_1_43; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10421 = _T_10420 | _T_10210; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_10212 = _T_4944 & ic_tag_valid_out_1_44; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10422 = _T_10421 | _T_10212; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_10214 = _T_4945 & ic_tag_valid_out_1_45; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10423 = _T_10422 | _T_10214; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_10216 = _T_4946 & ic_tag_valid_out_1_46; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10424 = _T_10423 | _T_10216; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_10218 = _T_4947 & ic_tag_valid_out_1_47; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10425 = _T_10424 | _T_10218; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_10220 = _T_4948 & ic_tag_valid_out_1_48; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10426 = _T_10425 | _T_10220; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_10222 = _T_4949 & ic_tag_valid_out_1_49; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10427 = _T_10426 | _T_10222; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_10224 = _T_4950 & ic_tag_valid_out_1_50; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10428 = _T_10427 | _T_10224; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_10226 = _T_4951 & ic_tag_valid_out_1_51; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10429 = _T_10428 | _T_10226; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_10228 = _T_4952 & ic_tag_valid_out_1_52; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10430 = _T_10429 | _T_10228; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_10230 = _T_4953 & ic_tag_valid_out_1_53; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10431 = _T_10430 | _T_10230; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_10232 = _T_4954 & ic_tag_valid_out_1_54; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10432 = _T_10431 | _T_10232; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_10234 = _T_4955 & ic_tag_valid_out_1_55; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10433 = _T_10432 | _T_10234; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_10236 = _T_4956 & ic_tag_valid_out_1_56; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10434 = _T_10433 | _T_10236; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_10238 = _T_4957 & ic_tag_valid_out_1_57; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10435 = _T_10434 | _T_10238; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_10240 = _T_4958 & ic_tag_valid_out_1_58; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10436 = _T_10435 | _T_10240; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_10242 = _T_4959 & ic_tag_valid_out_1_59; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10437 = _T_10436 | _T_10242; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_10244 = _T_4960 & ic_tag_valid_out_1_60; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10438 = _T_10437 | _T_10244; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_10246 = _T_4961 & ic_tag_valid_out_1_61; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10439 = _T_10438 | _T_10246; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_10248 = _T_4962 & ic_tag_valid_out_1_62; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10440 = _T_10439 | _T_10248; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_10250 = _T_4963 & ic_tag_valid_out_1_63; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10441 = _T_10440 | _T_10250; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_10252 = _T_4964 & ic_tag_valid_out_1_64; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10442 = _T_10441 | _T_10252; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_10254 = _T_4965 & ic_tag_valid_out_1_65; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10443 = _T_10442 | _T_10254; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_10256 = _T_4966 & ic_tag_valid_out_1_66; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10444 = _T_10443 | _T_10256; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_10258 = _T_4967 & ic_tag_valid_out_1_67; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10445 = _T_10444 | _T_10258; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_10260 = _T_4968 & ic_tag_valid_out_1_68; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10446 = _T_10445 | _T_10260; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_10262 = _T_4969 & ic_tag_valid_out_1_69; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10447 = _T_10446 | _T_10262; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_10264 = _T_4970 & ic_tag_valid_out_1_70; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10448 = _T_10447 | _T_10264; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_10266 = _T_4971 & ic_tag_valid_out_1_71; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10449 = _T_10448 | _T_10266; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_10268 = _T_4972 & ic_tag_valid_out_1_72; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10450 = _T_10449 | _T_10268; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_10270 = _T_4973 & ic_tag_valid_out_1_73; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10451 = _T_10450 | _T_10270; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_10272 = _T_4974 & ic_tag_valid_out_1_74; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10452 = _T_10451 | _T_10272; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_10274 = _T_4975 & ic_tag_valid_out_1_75; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10453 = _T_10452 | _T_10274; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_10276 = _T_4976 & ic_tag_valid_out_1_76; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10454 = _T_10453 | _T_10276; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_10278 = _T_4977 & ic_tag_valid_out_1_77; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10455 = _T_10454 | _T_10278; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_10280 = _T_4978 & ic_tag_valid_out_1_78; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10456 = _T_10455 | _T_10280; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_10282 = _T_4979 & ic_tag_valid_out_1_79; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10457 = _T_10456 | _T_10282; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_10284 = _T_4980 & ic_tag_valid_out_1_80; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10458 = _T_10457 | _T_10284; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_10286 = _T_4981 & ic_tag_valid_out_1_81; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10459 = _T_10458 | _T_10286; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_10288 = _T_4982 & ic_tag_valid_out_1_82; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10460 = _T_10459 | _T_10288; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_10290 = _T_4983 & ic_tag_valid_out_1_83; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10461 = _T_10460 | _T_10290; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_10292 = _T_4984 & ic_tag_valid_out_1_84; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10462 = _T_10461 | _T_10292; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_10294 = _T_4985 & ic_tag_valid_out_1_85; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10463 = _T_10462 | _T_10294; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_10296 = _T_4986 & ic_tag_valid_out_1_86; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10464 = _T_10463 | _T_10296; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_10298 = _T_4987 & ic_tag_valid_out_1_87; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10465 = _T_10464 | _T_10298; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_10300 = _T_4988 & ic_tag_valid_out_1_88; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10466 = _T_10465 | _T_10300; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_10302 = _T_4989 & ic_tag_valid_out_1_89; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10467 = _T_10466 | _T_10302; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_10304 = _T_4990 & ic_tag_valid_out_1_90; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10468 = _T_10467 | _T_10304; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_10306 = _T_4991 & ic_tag_valid_out_1_91; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10469 = _T_10468 | _T_10306; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_10308 = _T_4992 & ic_tag_valid_out_1_92; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10470 = _T_10469 | _T_10308; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_10310 = _T_4993 & ic_tag_valid_out_1_93; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10471 = _T_10470 | _T_10310; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_10312 = _T_4994 & ic_tag_valid_out_1_94; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10472 = _T_10471 | _T_10312; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_10314 = _T_4995 & ic_tag_valid_out_1_95; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10473 = _T_10472 | _T_10314; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_10316 = _T_4996 & ic_tag_valid_out_1_96; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10474 = _T_10473 | _T_10316; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_10318 = _T_4997 & ic_tag_valid_out_1_97; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10475 = _T_10474 | _T_10318; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_10320 = _T_4998 & ic_tag_valid_out_1_98; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10476 = _T_10475 | _T_10320; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_10322 = _T_4999 & ic_tag_valid_out_1_99; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10477 = _T_10476 | _T_10322; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_10324 = _T_5000 & ic_tag_valid_out_1_100; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10478 = _T_10477 | _T_10324; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_10326 = _T_5001 & ic_tag_valid_out_1_101; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10479 = _T_10478 | _T_10326; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_10328 = _T_5002 & ic_tag_valid_out_1_102; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10480 = _T_10479 | _T_10328; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_10330 = _T_5003 & ic_tag_valid_out_1_103; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10481 = _T_10480 | _T_10330; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_10332 = _T_5004 & ic_tag_valid_out_1_104; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10482 = _T_10481 | _T_10332; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_10334 = _T_5005 & ic_tag_valid_out_1_105; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10483 = _T_10482 | _T_10334; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_10336 = _T_5006 & ic_tag_valid_out_1_106; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10484 = _T_10483 | _T_10336; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_10338 = _T_5007 & ic_tag_valid_out_1_107; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10485 = _T_10484 | _T_10338; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_10340 = _T_5008 & ic_tag_valid_out_1_108; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10486 = _T_10485 | _T_10340; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_10342 = _T_5009 & ic_tag_valid_out_1_109; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10487 = _T_10486 | _T_10342; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_10344 = _T_5010 & ic_tag_valid_out_1_110; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10488 = _T_10487 | _T_10344; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_10346 = _T_5011 & ic_tag_valid_out_1_111; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10489 = _T_10488 | _T_10346; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_10348 = _T_5012 & ic_tag_valid_out_1_112; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10490 = _T_10489 | _T_10348; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_10350 = _T_5013 & ic_tag_valid_out_1_113; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10491 = _T_10490 | _T_10350; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_10352 = _T_5014 & ic_tag_valid_out_1_114; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10492 = _T_10491 | _T_10352; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_10354 = _T_5015 & ic_tag_valid_out_1_115; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10493 = _T_10492 | _T_10354; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_10356 = _T_5016 & ic_tag_valid_out_1_116; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10494 = _T_10493 | _T_10356; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_10358 = _T_5017 & ic_tag_valid_out_1_117; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10495 = _T_10494 | _T_10358; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_10360 = _T_5018 & ic_tag_valid_out_1_118; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10496 = _T_10495 | _T_10360; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_10362 = _T_5019 & ic_tag_valid_out_1_119; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10497 = _T_10496 | _T_10362; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_10364 = _T_5020 & ic_tag_valid_out_1_120; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10498 = _T_10497 | _T_10364; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_10366 = _T_5021 & ic_tag_valid_out_1_121; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10499 = _T_10498 | _T_10366; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_10368 = _T_5022 & ic_tag_valid_out_1_122; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10500 = _T_10499 | _T_10368; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_10370 = _T_5023 & ic_tag_valid_out_1_123; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10501 = _T_10500 | _T_10370; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_10372 = _T_5024 & ic_tag_valid_out_1_124; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10502 = _T_10501 | _T_10372; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_10374 = _T_5025 & ic_tag_valid_out_1_125; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10503 = _T_10502 | _T_10374; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_10376 = _T_5026 & ic_tag_valid_out_1_126; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10504 = _T_10503 | _T_10376; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_10378 = _T_5027 & ic_tag_valid_out_1_127; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10505 = _T_10504 | _T_10378; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_9741 = _T_4900 & ic_tag_valid_out_0_0; // @[ifu_mem_ctl.scala 656:8]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_9743 = _T_4901 & ic_tag_valid_out_0_1; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_9996 = _T_9741 | _T_9743; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_9745 = _T_4902 & ic_tag_valid_out_0_2; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_9997 = _T_9996 | _T_9745; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_9747 = _T_4903 & ic_tag_valid_out_0_3; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_9998 = _T_9997 | _T_9747; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_9749 = _T_4904 & ic_tag_valid_out_0_4; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_9999 = _T_9998 | _T_9749; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9751 = _T_4905 & ic_tag_valid_out_0_5; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10000 = _T_9999 | _T_9751; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9753 = _T_4906 & ic_tag_valid_out_0_6; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10001 = _T_10000 | _T_9753; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9755 = _T_4907 & ic_tag_valid_out_0_7; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10002 = _T_10001 | _T_9755; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9757 = _T_4908 & ic_tag_valid_out_0_8; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10003 = _T_10002 | _T_9757; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9759 = _T_4909 & ic_tag_valid_out_0_9; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10004 = _T_10003 | _T_9759; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9761 = _T_4910 & ic_tag_valid_out_0_10; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10005 = _T_10004 | _T_9761; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9763 = _T_4911 & ic_tag_valid_out_0_11; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10006 = _T_10005 | _T_9763; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9765 = _T_4912 & ic_tag_valid_out_0_12; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10007 = _T_10006 | _T_9765; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9767 = _T_4913 & ic_tag_valid_out_0_13; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10008 = _T_10007 | _T_9767; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9769 = _T_4914 & ic_tag_valid_out_0_14; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10009 = _T_10008 | _T_9769; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9771 = _T_4915 & ic_tag_valid_out_0_15; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10010 = _T_10009 | _T_9771; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9773 = _T_4916 & ic_tag_valid_out_0_16; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10011 = _T_10010 | _T_9773; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9775 = _T_4917 & ic_tag_valid_out_0_17; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10012 = _T_10011 | _T_9775; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9777 = _T_4918 & ic_tag_valid_out_0_18; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10013 = _T_10012 | _T_9777; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9779 = _T_4919 & ic_tag_valid_out_0_19; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10014 = _T_10013 | _T_9779; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9781 = _T_4920 & ic_tag_valid_out_0_20; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10015 = _T_10014 | _T_9781; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9783 = _T_4921 & ic_tag_valid_out_0_21; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10016 = _T_10015 | _T_9783; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9785 = _T_4922 & ic_tag_valid_out_0_22; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10017 = _T_10016 | _T_9785; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9787 = _T_4923 & ic_tag_valid_out_0_23; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10018 = _T_10017 | _T_9787; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9789 = _T_4924 & ic_tag_valid_out_0_24; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10019 = _T_10018 | _T_9789; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9791 = _T_4925 & ic_tag_valid_out_0_25; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10020 = _T_10019 | _T_9791; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9793 = _T_4926 & ic_tag_valid_out_0_26; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10021 = _T_10020 | _T_9793; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9795 = _T_4927 & ic_tag_valid_out_0_27; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10022 = _T_10021 | _T_9795; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9797 = _T_4928 & ic_tag_valid_out_0_28; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10023 = _T_10022 | _T_9797; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9799 = _T_4929 & ic_tag_valid_out_0_29; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10024 = _T_10023 | _T_9799; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9801 = _T_4930 & ic_tag_valid_out_0_30; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10025 = _T_10024 | _T_9801; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9803 = _T_4931 & ic_tag_valid_out_0_31; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10026 = _T_10025 | _T_9803; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9805 = _T_4932 & ic_tag_valid_out_0_32; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10027 = _T_10026 | _T_9805; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9807 = _T_4933 & ic_tag_valid_out_0_33; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10028 = _T_10027 | _T_9807; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9809 = _T_4934 & ic_tag_valid_out_0_34; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10029 = _T_10028 | _T_9809; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9811 = _T_4935 & ic_tag_valid_out_0_35; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10030 = _T_10029 | _T_9811; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9813 = _T_4936 & ic_tag_valid_out_0_36; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10031 = _T_10030 | _T_9813; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9815 = _T_4937 & ic_tag_valid_out_0_37; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10032 = _T_10031 | _T_9815; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9817 = _T_4938 & ic_tag_valid_out_0_38; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10033 = _T_10032 | _T_9817; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9819 = _T_4939 & ic_tag_valid_out_0_39; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10034 = _T_10033 | _T_9819; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9821 = _T_4940 & ic_tag_valid_out_0_40; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10035 = _T_10034 | _T_9821; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9823 = _T_4941 & ic_tag_valid_out_0_41; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10036 = _T_10035 | _T_9823; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9825 = _T_4942 & ic_tag_valid_out_0_42; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10037 = _T_10036 | _T_9825; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9827 = _T_4943 & ic_tag_valid_out_0_43; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10038 = _T_10037 | _T_9827; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9829 = _T_4944 & ic_tag_valid_out_0_44; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10039 = _T_10038 | _T_9829; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9831 = _T_4945 & ic_tag_valid_out_0_45; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10040 = _T_10039 | _T_9831; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9833 = _T_4946 & ic_tag_valid_out_0_46; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10041 = _T_10040 | _T_9833; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9835 = _T_4947 & ic_tag_valid_out_0_47; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10042 = _T_10041 | _T_9835; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9837 = _T_4948 & ic_tag_valid_out_0_48; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10043 = _T_10042 | _T_9837; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9839 = _T_4949 & ic_tag_valid_out_0_49; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10044 = _T_10043 | _T_9839; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9841 = _T_4950 & ic_tag_valid_out_0_50; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10045 = _T_10044 | _T_9841; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9843 = _T_4951 & ic_tag_valid_out_0_51; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10046 = _T_10045 | _T_9843; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9845 = _T_4952 & ic_tag_valid_out_0_52; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10047 = _T_10046 | _T_9845; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9847 = _T_4953 & ic_tag_valid_out_0_53; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10048 = _T_10047 | _T_9847; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9849 = _T_4954 & ic_tag_valid_out_0_54; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10049 = _T_10048 | _T_9849; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9851 = _T_4955 & ic_tag_valid_out_0_55; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10050 = _T_10049 | _T_9851; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9853 = _T_4956 & ic_tag_valid_out_0_56; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10051 = _T_10050 | _T_9853; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9855 = _T_4957 & ic_tag_valid_out_0_57; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10052 = _T_10051 | _T_9855; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9857 = _T_4958 & ic_tag_valid_out_0_58; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10053 = _T_10052 | _T_9857; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9859 = _T_4959 & ic_tag_valid_out_0_59; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10054 = _T_10053 | _T_9859; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9861 = _T_4960 & ic_tag_valid_out_0_60; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10055 = _T_10054 | _T_9861; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9863 = _T_4961 & ic_tag_valid_out_0_61; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10056 = _T_10055 | _T_9863; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9865 = _T_4962 & ic_tag_valid_out_0_62; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10057 = _T_10056 | _T_9865; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9867 = _T_4963 & ic_tag_valid_out_0_63; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10058 = _T_10057 | _T_9867; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9869 = _T_4964 & ic_tag_valid_out_0_64; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10059 = _T_10058 | _T_9869; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9871 = _T_4965 & ic_tag_valid_out_0_65; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10060 = _T_10059 | _T_9871; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9873 = _T_4966 & ic_tag_valid_out_0_66; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10061 = _T_10060 | _T_9873; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9875 = _T_4967 & ic_tag_valid_out_0_67; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10062 = _T_10061 | _T_9875; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9877 = _T_4968 & ic_tag_valid_out_0_68; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10063 = _T_10062 | _T_9877; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9879 = _T_4969 & ic_tag_valid_out_0_69; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10064 = _T_10063 | _T_9879; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9881 = _T_4970 & ic_tag_valid_out_0_70; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10065 = _T_10064 | _T_9881; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9883 = _T_4971 & ic_tag_valid_out_0_71; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10066 = _T_10065 | _T_9883; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9885 = _T_4972 & ic_tag_valid_out_0_72; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10067 = _T_10066 | _T_9885; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9887 = _T_4973 & ic_tag_valid_out_0_73; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10068 = _T_10067 | _T_9887; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9889 = _T_4974 & ic_tag_valid_out_0_74; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10069 = _T_10068 | _T_9889; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9891 = _T_4975 & ic_tag_valid_out_0_75; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10070 = _T_10069 | _T_9891; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9893 = _T_4976 & ic_tag_valid_out_0_76; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10071 = _T_10070 | _T_9893; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9895 = _T_4977 & ic_tag_valid_out_0_77; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10072 = _T_10071 | _T_9895; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9897 = _T_4978 & ic_tag_valid_out_0_78; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10073 = _T_10072 | _T_9897; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9899 = _T_4979 & ic_tag_valid_out_0_79; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10074 = _T_10073 | _T_9899; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9901 = _T_4980 & ic_tag_valid_out_0_80; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10075 = _T_10074 | _T_9901; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9903 = _T_4981 & ic_tag_valid_out_0_81; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10076 = _T_10075 | _T_9903; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9905 = _T_4982 & ic_tag_valid_out_0_82; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10077 = _T_10076 | _T_9905; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9907 = _T_4983 & ic_tag_valid_out_0_83; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10078 = _T_10077 | _T_9907; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9909 = _T_4984 & ic_tag_valid_out_0_84; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10079 = _T_10078 | _T_9909; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9911 = _T_4985 & ic_tag_valid_out_0_85; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10080 = _T_10079 | _T_9911; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9913 = _T_4986 & ic_tag_valid_out_0_86; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10081 = _T_10080 | _T_9913; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9915 = _T_4987 & ic_tag_valid_out_0_87; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10082 = _T_10081 | _T_9915; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9917 = _T_4988 & ic_tag_valid_out_0_88; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10083 = _T_10082 | _T_9917; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9919 = _T_4989 & ic_tag_valid_out_0_89; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10084 = _T_10083 | _T_9919; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9921 = _T_4990 & ic_tag_valid_out_0_90; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10085 = _T_10084 | _T_9921; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9923 = _T_4991 & ic_tag_valid_out_0_91; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10086 = _T_10085 | _T_9923; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9925 = _T_4992 & ic_tag_valid_out_0_92; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10087 = _T_10086 | _T_9925; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9927 = _T_4993 & ic_tag_valid_out_0_93; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10088 = _T_10087 | _T_9927; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9929 = _T_4994 & ic_tag_valid_out_0_94; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10089 = _T_10088 | _T_9929; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9931 = _T_4995 & ic_tag_valid_out_0_95; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10090 = _T_10089 | _T_9931; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9933 = _T_4996 & ic_tag_valid_out_0_96; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10091 = _T_10090 | _T_9933; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9935 = _T_4997 & ic_tag_valid_out_0_97; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10092 = _T_10091 | _T_9935; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9937 = _T_4998 & ic_tag_valid_out_0_98; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10093 = _T_10092 | _T_9937; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9939 = _T_4999 & ic_tag_valid_out_0_99; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10094 = _T_10093 | _T_9939; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9941 = _T_5000 & ic_tag_valid_out_0_100; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10095 = _T_10094 | _T_9941; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9943 = _T_5001 & ic_tag_valid_out_0_101; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10096 = _T_10095 | _T_9943; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9945 = _T_5002 & ic_tag_valid_out_0_102; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10097 = _T_10096 | _T_9945; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9947 = _T_5003 & ic_tag_valid_out_0_103; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10098 = _T_10097 | _T_9947; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9949 = _T_5004 & ic_tag_valid_out_0_104; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10099 = _T_10098 | _T_9949; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9951 = _T_5005 & ic_tag_valid_out_0_105; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10100 = _T_10099 | _T_9951; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9953 = _T_5006 & ic_tag_valid_out_0_106; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10101 = _T_10100 | _T_9953; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9955 = _T_5007 & ic_tag_valid_out_0_107; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10102 = _T_10101 | _T_9955; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9957 = _T_5008 & ic_tag_valid_out_0_108; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10103 = _T_10102 | _T_9957; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9959 = _T_5009 & ic_tag_valid_out_0_109; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10104 = _T_10103 | _T_9959; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9961 = _T_5010 & ic_tag_valid_out_0_110; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10105 = _T_10104 | _T_9961; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9963 = _T_5011 & ic_tag_valid_out_0_111; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10106 = _T_10105 | _T_9963; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9965 = _T_5012 & ic_tag_valid_out_0_112; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10107 = _T_10106 | _T_9965; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9967 = _T_5013 & ic_tag_valid_out_0_113; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10108 = _T_10107 | _T_9967; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9969 = _T_5014 & ic_tag_valid_out_0_114; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10109 = _T_10108 | _T_9969; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9971 = _T_5015 & ic_tag_valid_out_0_115; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10110 = _T_10109 | _T_9971; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9973 = _T_5016 & ic_tag_valid_out_0_116; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10111 = _T_10110 | _T_9973; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9975 = _T_5017 & ic_tag_valid_out_0_117; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10112 = _T_10111 | _T_9975; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9977 = _T_5018 & ic_tag_valid_out_0_118; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10113 = _T_10112 | _T_9977; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9979 = _T_5019 & ic_tag_valid_out_0_119; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10114 = _T_10113 | _T_9979; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9981 = _T_5020 & ic_tag_valid_out_0_120; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10115 = _T_10114 | _T_9981; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9983 = _T_5021 & ic_tag_valid_out_0_121; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10116 = _T_10115 | _T_9983; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9985 = _T_5022 & ic_tag_valid_out_0_122; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10117 = _T_10116 | _T_9985; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9987 = _T_5023 & ic_tag_valid_out_0_123; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10118 = _T_10117 | _T_9987; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9989 = _T_5024 & ic_tag_valid_out_0_124; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10119 = _T_10118 | _T_9989; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9991 = _T_5025 & ic_tag_valid_out_0_125; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10120 = _T_10119 | _T_9991; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9993 = _T_5026 & ic_tag_valid_out_0_126; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10121 = _T_10120 | _T_9993; // @[ifu_mem_ctl.scala 656:85]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9995 = _T_5027 & ic_tag_valid_out_0_127; // @[ifu_mem_ctl.scala 656:8]
  wire  _T_10122 = _T_10121 | _T_9995; // @[ifu_mem_ctl.scala 656:85]
  wire [1:0] ic_tag_valid_unq = {_T_10505,_T_10122}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[Reg.scala 27:20]
  wire [1:0] _T_10545 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10546 = ic_debug_way_ff & _T_10545; // @[ifu_mem_ctl.scala 705:67]
  wire [1:0] _T_10547 = ic_tag_valid_unq & _T_10546; // @[ifu_mem_ctl.scala 705:48]
  wire  ic_debug_tag_val_rd_out = |_T_10547; // @[ifu_mem_ctl.scala 705:115]
  wire [70:0] _T_1236 = {2'h0,io_ic_tag_debug_rd_data[25:21],32'h0,io_ic_tag_debug_rd_data[20:0],6'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1237; // @[Reg.scala 27:20]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2657; // @[ifu_mem_ctl.scala 270:84]
  wire  _T_1271 = ifu_wr_cumulative_err ^ ifu_wr_data_comb_err_ff; // @[lib.scala 453:21]
  wire  _T_1272 = |_T_1271; // @[lib.scala 453:29]
  wire  _T_1287 = _T_1280 | fetch_req_iccm_f; // @[ifu_mem_ctl.scala 280:61]
  wire  _T_1288 = _T_1287 | sel_ic_data; // @[ifu_mem_ctl.scala 280:80]
  wire [63:0] _T_1290 = _T_1288 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] ic_final_data = _T_1290 & io_ic_rd_data; // @[ifu_mem_ctl.scala 280:95]
  wire [63:0] _T_1292 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1293 = _T_1292 & io_iccm_rd_data; // @[ifu_mem_ctl.scala 284:72]
  wire [63:0] _T_1295 = _T_1280 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2153 = ~ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 350:31]
  wire  _T_1666 = ~ifu_fetch_addr_int_f[1]; // @[ifu_mem_ctl.scala 346:38]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1667 = byp_fetch_index_inc_0 == 4'h0; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1715 = _T_1667 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1670 = byp_fetch_index_inc_0 == 4'h1; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1716 = _T_1670 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1731 = _T_1715 | _T_1716; // @[Mux.scala 27:72]
  wire  _T_1673 = byp_fetch_index_inc_0 == 4'h2; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1717 = _T_1673 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1732 = _T_1731 | _T_1717; // @[Mux.scala 27:72]
  wire  _T_1676 = byp_fetch_index_inc_0 == 4'h3; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1718 = _T_1676 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1733 = _T_1732 | _T_1718; // @[Mux.scala 27:72]
  wire  _T_1679 = byp_fetch_index_inc_0 == 4'h4; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1719 = _T_1679 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1734 = _T_1733 | _T_1719; // @[Mux.scala 27:72]
  wire  _T_1682 = byp_fetch_index_inc_0 == 4'h5; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1720 = _T_1682 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1735 = _T_1734 | _T_1720; // @[Mux.scala 27:72]
  wire  _T_1685 = byp_fetch_index_inc_0 == 4'h6; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1721 = _T_1685 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1736 = _T_1735 | _T_1721; // @[Mux.scala 27:72]
  wire  _T_1688 = byp_fetch_index_inc_0 == 4'h7; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1722 = _T_1688 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1737 = _T_1736 | _T_1722; // @[Mux.scala 27:72]
  wire  _T_1691 = byp_fetch_index_inc_0 == 4'h8; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1723 = _T_1691 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1738 = _T_1737 | _T_1723; // @[Mux.scala 27:72]
  wire  _T_1694 = byp_fetch_index_inc_0 == 4'h9; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1724 = _T_1694 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1739 = _T_1738 | _T_1724; // @[Mux.scala 27:72]
  wire  _T_1697 = byp_fetch_index_inc_0 == 4'ha; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1725 = _T_1697 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1740 = _T_1739 | _T_1725; // @[Mux.scala 27:72]
  wire  _T_1700 = byp_fetch_index_inc_0 == 4'hb; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1726 = _T_1700 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1741 = _T_1740 | _T_1726; // @[Mux.scala 27:72]
  wire  _T_1703 = byp_fetch_index_inc_0 == 4'hc; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1727 = _T_1703 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1742 = _T_1741 | _T_1727; // @[Mux.scala 27:72]
  wire  _T_1706 = byp_fetch_index_inc_0 == 4'hd; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1728 = _T_1706 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1743 = _T_1742 | _T_1728; // @[Mux.scala 27:72]
  wire  _T_1709 = byp_fetch_index_inc_0 == 4'he; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1729 = _T_1709 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1744 = _T_1743 | _T_1729; // @[Mux.scala 27:72]
  wire  _T_1712 = byp_fetch_index_inc_0 == 4'hf; // @[ifu_mem_ctl.scala 347:73]
  wire [15:0] _T_1730 = _T_1712 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1745 = _T_1744 | _T_1730; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1747 = byp_fetch_index_1 == 4'h0; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1795 = _T_1747 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1750 = byp_fetch_index_1 == 4'h1; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1796 = _T_1750 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1811 = _T_1795 | _T_1796; // @[Mux.scala 27:72]
  wire  _T_1753 = byp_fetch_index_1 == 4'h2; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1797 = _T_1753 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1812 = _T_1811 | _T_1797; // @[Mux.scala 27:72]
  wire  _T_1756 = byp_fetch_index_1 == 4'h3; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1798 = _T_1756 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1813 = _T_1812 | _T_1798; // @[Mux.scala 27:72]
  wire  _T_1759 = byp_fetch_index_1 == 4'h4; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1799 = _T_1759 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1814 = _T_1813 | _T_1799; // @[Mux.scala 27:72]
  wire  _T_1762 = byp_fetch_index_1 == 4'h5; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1800 = _T_1762 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1815 = _T_1814 | _T_1800; // @[Mux.scala 27:72]
  wire  _T_1765 = byp_fetch_index_1 == 4'h6; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1801 = _T_1765 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1816 = _T_1815 | _T_1801; // @[Mux.scala 27:72]
  wire  _T_1768 = byp_fetch_index_1 == 4'h7; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1802 = _T_1768 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1817 = _T_1816 | _T_1802; // @[Mux.scala 27:72]
  wire  _T_1771 = byp_fetch_index_1 == 4'h8; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1803 = _T_1771 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1818 = _T_1817 | _T_1803; // @[Mux.scala 27:72]
  wire  _T_1774 = byp_fetch_index_1 == 4'h9; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1804 = _T_1774 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1819 = _T_1818 | _T_1804; // @[Mux.scala 27:72]
  wire  _T_1777 = byp_fetch_index_1 == 4'ha; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1805 = _T_1777 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1820 = _T_1819 | _T_1805; // @[Mux.scala 27:72]
  wire  _T_1780 = byp_fetch_index_1 == 4'hb; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1806 = _T_1780 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1821 = _T_1820 | _T_1806; // @[Mux.scala 27:72]
  wire  _T_1783 = byp_fetch_index_1 == 4'hc; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1807 = _T_1783 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1822 = _T_1821 | _T_1807; // @[Mux.scala 27:72]
  wire  _T_1786 = byp_fetch_index_1 == 4'hd; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1808 = _T_1786 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1823 = _T_1822 | _T_1808; // @[Mux.scala 27:72]
  wire  _T_1789 = byp_fetch_index_1 == 4'he; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1809 = _T_1789 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1824 = _T_1823 | _T_1809; // @[Mux.scala 27:72]
  wire  _T_1792 = byp_fetch_index_1 == 4'hf; // @[ifu_mem_ctl.scala 347:179]
  wire [31:0] _T_1810 = _T_1792 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1825 = _T_1824 | _T_1810; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1827 = byp_fetch_index_0 == 4'h0; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1875 = _T_1827 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1830 = byp_fetch_index_0 == 4'h1; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1876 = _T_1830 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1891 = _T_1875 | _T_1876; // @[Mux.scala 27:72]
  wire  _T_1833 = byp_fetch_index_0 == 4'h2; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1877 = _T_1833 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1892 = _T_1891 | _T_1877; // @[Mux.scala 27:72]
  wire  _T_1836 = byp_fetch_index_0 == 4'h3; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1878 = _T_1836 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1893 = _T_1892 | _T_1878; // @[Mux.scala 27:72]
  wire  _T_1839 = byp_fetch_index_0 == 4'h4; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1879 = _T_1839 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1894 = _T_1893 | _T_1879; // @[Mux.scala 27:72]
  wire  _T_1842 = byp_fetch_index_0 == 4'h5; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1880 = _T_1842 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1895 = _T_1894 | _T_1880; // @[Mux.scala 27:72]
  wire  _T_1845 = byp_fetch_index_0 == 4'h6; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1881 = _T_1845 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1896 = _T_1895 | _T_1881; // @[Mux.scala 27:72]
  wire  _T_1848 = byp_fetch_index_0 == 4'h7; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1882 = _T_1848 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1897 = _T_1896 | _T_1882; // @[Mux.scala 27:72]
  wire  _T_1851 = byp_fetch_index_0 == 4'h8; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1883 = _T_1851 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1898 = _T_1897 | _T_1883; // @[Mux.scala 27:72]
  wire  _T_1854 = byp_fetch_index_0 == 4'h9; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1884 = _T_1854 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1899 = _T_1898 | _T_1884; // @[Mux.scala 27:72]
  wire  _T_1857 = byp_fetch_index_0 == 4'ha; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1885 = _T_1857 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1900 = _T_1899 | _T_1885; // @[Mux.scala 27:72]
  wire  _T_1860 = byp_fetch_index_0 == 4'hb; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1886 = _T_1860 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1901 = _T_1900 | _T_1886; // @[Mux.scala 27:72]
  wire  _T_1863 = byp_fetch_index_0 == 4'hc; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1887 = _T_1863 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1902 = _T_1901 | _T_1887; // @[Mux.scala 27:72]
  wire  _T_1866 = byp_fetch_index_0 == 4'hd; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1888 = _T_1866 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1903 = _T_1902 | _T_1888; // @[Mux.scala 27:72]
  wire  _T_1869 = byp_fetch_index_0 == 4'he; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1889 = _T_1869 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1904 = _T_1903 | _T_1889; // @[Mux.scala 27:72]
  wire  _T_1872 = byp_fetch_index_0 == 4'hf; // @[ifu_mem_ctl.scala 347:285]
  wire [31:0] _T_1890 = _T_1872 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1905 = _T_1904 | _T_1890; // @[Mux.scala 27:72]
  wire [79:0] _T_1908 = {_T_1745,_T_1825,_T_1905}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1909 = byp_fetch_index_inc_1 == 4'h0; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1957 = _T_1909 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1912 = byp_fetch_index_inc_1 == 4'h1; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1958 = _T_1912 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1973 = _T_1957 | _T_1958; // @[Mux.scala 27:72]
  wire  _T_1915 = byp_fetch_index_inc_1 == 4'h2; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1959 = _T_1915 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1974 = _T_1973 | _T_1959; // @[Mux.scala 27:72]
  wire  _T_1918 = byp_fetch_index_inc_1 == 4'h3; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1960 = _T_1918 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1975 = _T_1974 | _T_1960; // @[Mux.scala 27:72]
  wire  _T_1921 = byp_fetch_index_inc_1 == 4'h4; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1961 = _T_1921 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1976 = _T_1975 | _T_1961; // @[Mux.scala 27:72]
  wire  _T_1924 = byp_fetch_index_inc_1 == 4'h5; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1962 = _T_1924 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1977 = _T_1976 | _T_1962; // @[Mux.scala 27:72]
  wire  _T_1927 = byp_fetch_index_inc_1 == 4'h6; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1963 = _T_1927 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1978 = _T_1977 | _T_1963; // @[Mux.scala 27:72]
  wire  _T_1930 = byp_fetch_index_inc_1 == 4'h7; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1964 = _T_1930 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1979 = _T_1978 | _T_1964; // @[Mux.scala 27:72]
  wire  _T_1933 = byp_fetch_index_inc_1 == 4'h8; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1965 = _T_1933 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1980 = _T_1979 | _T_1965; // @[Mux.scala 27:72]
  wire  _T_1936 = byp_fetch_index_inc_1 == 4'h9; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1966 = _T_1936 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1981 = _T_1980 | _T_1966; // @[Mux.scala 27:72]
  wire  _T_1939 = byp_fetch_index_inc_1 == 4'ha; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1967 = _T_1939 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1982 = _T_1981 | _T_1967; // @[Mux.scala 27:72]
  wire  _T_1942 = byp_fetch_index_inc_1 == 4'hb; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1968 = _T_1942 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1983 = _T_1982 | _T_1968; // @[Mux.scala 27:72]
  wire  _T_1945 = byp_fetch_index_inc_1 == 4'hc; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1969 = _T_1945 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1984 = _T_1983 | _T_1969; // @[Mux.scala 27:72]
  wire  _T_1948 = byp_fetch_index_inc_1 == 4'hd; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1970 = _T_1948 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1985 = _T_1984 | _T_1970; // @[Mux.scala 27:72]
  wire  _T_1951 = byp_fetch_index_inc_1 == 4'he; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1971 = _T_1951 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1986 = _T_1985 | _T_1971; // @[Mux.scala 27:72]
  wire  _T_1954 = byp_fetch_index_inc_1 == 4'hf; // @[ifu_mem_ctl.scala 348:73]
  wire [15:0] _T_1972 = _T_1954 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1987 = _T_1986 | _T_1972; // @[Mux.scala 27:72]
  wire [31:0] _T_2037 = _T_1667 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2038 = _T_1670 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2053 = _T_2037 | _T_2038; // @[Mux.scala 27:72]
  wire [31:0] _T_2039 = _T_1673 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2054 = _T_2053 | _T_2039; // @[Mux.scala 27:72]
  wire [31:0] _T_2040 = _T_1676 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2055 = _T_2054 | _T_2040; // @[Mux.scala 27:72]
  wire [31:0] _T_2041 = _T_1679 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2056 = _T_2055 | _T_2041; // @[Mux.scala 27:72]
  wire [31:0] _T_2042 = _T_1682 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2057 = _T_2056 | _T_2042; // @[Mux.scala 27:72]
  wire [31:0] _T_2043 = _T_1685 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2058 = _T_2057 | _T_2043; // @[Mux.scala 27:72]
  wire [31:0] _T_2044 = _T_1688 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2059 = _T_2058 | _T_2044; // @[Mux.scala 27:72]
  wire [31:0] _T_2045 = _T_1691 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2060 = _T_2059 | _T_2045; // @[Mux.scala 27:72]
  wire [31:0] _T_2046 = _T_1694 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2061 = _T_2060 | _T_2046; // @[Mux.scala 27:72]
  wire [31:0] _T_2047 = _T_1697 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2062 = _T_2061 | _T_2047; // @[Mux.scala 27:72]
  wire [31:0] _T_2048 = _T_1700 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2063 = _T_2062 | _T_2048; // @[Mux.scala 27:72]
  wire [31:0] _T_2049 = _T_1703 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2064 = _T_2063 | _T_2049; // @[Mux.scala 27:72]
  wire [31:0] _T_2050 = _T_1706 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2065 = _T_2064 | _T_2050; // @[Mux.scala 27:72]
  wire [31:0] _T_2051 = _T_1709 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2066 = _T_2065 | _T_2051; // @[Mux.scala 27:72]
  wire [31:0] _T_2052 = _T_1712 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2067 = _T_2066 | _T_2052; // @[Mux.scala 27:72]
  wire [79:0] _T_2150 = {_T_1987,_T_2067,_T_1825}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1666 ? _T_1908 : _T_2150; // @[ifu_mem_ctl.scala 346:37]
  wire [79:0] _T_2155 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2153 ? ic_byp_data_only_pre_new : _T_2155; // @[ifu_mem_ctl.scala 350:30]
  wire [79:0] _GEN_517 = {{16'd0}, _T_1295}; // @[ifu_mem_ctl.scala 284:117]
  wire [79:0] _T_1296 = _GEN_517 & ic_byp_data_only_new; // @[ifu_mem_ctl.scala 284:117]
  wire [79:0] _GEN_518 = {{16'd0}, _T_1293}; // @[ifu_mem_ctl.scala 284:91]
  wire [79:0] ic_premux_data_temp = _GEN_518 | _T_1296; // @[ifu_mem_ctl.scala 284:91]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_339; // @[ifu_mem_ctl.scala 291:38]
  wire [1:0] _T_1301 = ifc_region_acc_fault_final_f ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_1302 = _T_1301 | ifc_bus_acc_fault_f; // @[ifu_mem_ctl.scala 293:65]
  wire [1:0] _T_1305 = _T_339 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_1307 = |io_iccm_rd_ecc_double_err; // @[ifu_mem_ctl.scala 294:62]
  reg  ifc_region_acc_fault_memory_f; // @[Reg.scala 27:20]
  wire [1:0] _T_1309 = ifc_region_acc_fault_memory_f ? 2'h3 : 2'h0; // @[ifu_mem_ctl.scala 294:108]
  wire [1:0] _T_1310 = ifc_region_acc_fault_f ? 2'h2 : _T_1309; // @[ifu_mem_ctl.scala 294:75]
  wire  _T_1312 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[ifu_mem_ctl.scala 296:45]
  wire  _T_1314 = byp_fetch_index == 5'h1f; // @[ifu_mem_ctl.scala 296:80]
  wire  _T_1315 = ~_T_1314; // @[ifu_mem_ctl.scala 296:71]
  wire  _T_1316 = _T_1312 & _T_1315; // @[ifu_mem_ctl.scala 296:69]
  wire  _T_1317 = err_stop_state != 2'h2; // @[ifu_mem_ctl.scala 296:131]
  wire  _T_1318 = _T_1316 & _T_1317; // @[ifu_mem_ctl.scala 296:114]
  wire [6:0] _T_1390 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1}; // @[Cat.scala 29:58]
  wire  _T_1396 = ic_miss_buff_data_error[0] & _T_1362; // @[ifu_mem_ctl.scala 314:32]
  wire  _T_2734 = |io_ifu_axi_r_bits_resp; // @[ifu_mem_ctl.scala 521:54]
  wire  _T_2735 = _T_2734 & _T_16; // @[ifu_mem_ctl.scala 521:57]
  wire  bus_ifu_wr_data_error = _T_2735 & miss_pending; // @[ifu_mem_ctl.scala 521:75]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1396; // @[ifu_mem_ctl.scala 313:72]
  wire  _T_1400 = ic_miss_buff_data_error[1] & _T_1362; // @[ifu_mem_ctl.scala 314:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1400; // @[ifu_mem_ctl.scala 313:72]
  wire  _T_1404 = ic_miss_buff_data_error[2] & _T_1362; // @[ifu_mem_ctl.scala 314:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1404; // @[ifu_mem_ctl.scala 313:72]
  wire  _T_1408 = ic_miss_buff_data_error[3] & _T_1362; // @[ifu_mem_ctl.scala 314:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1408; // @[ifu_mem_ctl.scala 313:72]
  wire  _T_1412 = ic_miss_buff_data_error[4] & _T_1362; // @[ifu_mem_ctl.scala 314:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1412; // @[ifu_mem_ctl.scala 313:72]
  wire  _T_1416 = ic_miss_buff_data_error[5] & _T_1362; // @[ifu_mem_ctl.scala 314:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1416; // @[ifu_mem_ctl.scala 313:72]
  wire  _T_1420 = ic_miss_buff_data_error[6] & _T_1362; // @[ifu_mem_ctl.scala 314:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1420; // @[ifu_mem_ctl.scala 313:72]
  wire  _T_1424 = ic_miss_buff_data_error[7] & _T_1362; // @[ifu_mem_ctl.scala 314:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1424; // @[ifu_mem_ctl.scala 313:72]
  wire [6:0] _T_1430 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1}; // @[Cat.scala 29:58]
  wire  _T_1553 = ic_crit_wd_rdy_new_in ^ ic_crit_wd_rdy_new_ff; // @[lib.scala 453:21]
  wire  _T_1554 = |_T_1553; // @[lib.scala 453:29]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2521 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2529 = _T_9 & _T_339; // @[ifu_mem_ctl.scala 394:82]
  wire  _T_2530 = _T_2529 | io_iccm_dma_sb_error; // @[ifu_mem_ctl.scala 394:105]
  wire  _T_2532 = _T_2530 & _T_2653; // @[ifu_mem_ctl.scala 394:129]
  wire  _T_2533 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2534 = io_dec_tlu_flush_lower_wb | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 399:50]
  wire  _T_2536 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2543 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2545 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_60 = _T_2543 | _T_2545; // @[Conditional.scala 39:67]
  wire  _GEN_62 = _T_2536 ? _T_2534 : _GEN_60; // @[Conditional.scala 39:67]
  wire  _GEN_64 = _T_2533 ? _T_2534 : _GEN_62; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2521 ? _T_2532 : _GEN_64; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2521 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2535 = io_dec_tlu_flush_lower_wb & io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu_mem_ctl.scala 400:56]
  wire  _GEN_65 = _T_2533 & _T_2535; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2521 ? 1'h0 : _GEN_65; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[Reg.scala 27:20]
  wire  _T_2516 = _T_10 ^ dma_sb_err_state_ff; // @[lib.scala 475:21]
  wire  _T_2517 = |_T_2516; // @[lib.scala 475:29]
  wire  _T_2519 = ~dma_sb_err_state_ff; // @[ifu_mem_ctl.scala 385:49]
  wire  _T_2523 = io_dec_mem_ctrl_ifu_ic_error_start & _T_339; // @[ifu_mem_ctl.scala 393:104]
  wire  _T_2537 = ~io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu_mem_ctl.scala 403:30]
  wire  _T_2538 = _T_2537 & io_dec_tlu_flush_lower_wb; // @[ifu_mem_ctl.scala 403:68]
  wire  _T_2539 = _T_2538 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 403:98]
  wire  _T_2548 = perr_state == 3'h2; // @[ifu_mem_ctl.scala 423:79]
  wire  _T_2549 = io_dec_mem_ctrl_dec_tlu_flush_err_wb & _T_2548; // @[ifu_mem_ctl.scala 423:65]
  wire  _T_2551 = _T_2549 & _T_2653; // @[ifu_mem_ctl.scala 423:94]
  wire  _T_2553 = io_dec_tlu_flush_lower_wb | io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 426:59]
  wire  _T_2554 = _T_2553 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 426:99]
  wire  _T_2568 = _T_2553 | io_ifu_fetch_val[0]; // @[ifu_mem_ctl.scala 429:94]
  wire  _T_2569 = _T_2568 | ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 429:116]
  wire  _T_2570 = _T_2569 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 429:139]
  wire  _T_2590 = _T_2568 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 436:116]
  wire  _T_2598 = io_dec_tlu_flush_lower_wb & _T_2537; // @[ifu_mem_ctl.scala 441:60]
  wire  _T_2599 = _T_2598 | io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 441:101]
  wire  _T_2600 = _T_2599 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 441:141]
  wire  _GEN_72 = _T_2596 & _T_2554; // @[Conditional.scala 39:67]
  wire  _GEN_75 = _T_2579 ? _T_2590 : _GEN_72; // @[Conditional.scala 39:67]
  wire  _GEN_77 = _T_2579 | _T_2596; // @[Conditional.scala 39:67]
  wire  _GEN_79 = _T_2552 ? _T_2570 : _GEN_75; // @[Conditional.scala 39:67]
  wire  _GEN_81 = _T_2552 | _GEN_77; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2547 ? _T_2551 : _GEN_79; // @[Conditional.scala 40:58]
  wire  _T_2608 = io_ifu_bus_clk_en ^ bus_ifu_bus_clk_en_ff; // @[lib.scala 475:21]
  wire  _T_2609 = |_T_2608; // @[lib.scala 475:29]
  wire  _T_2612 = scnd_miss_req_in ^ scnd_miss_req_q; // @[lib.scala 475:21]
  wire  _T_2613 = |_T_2612; // @[lib.scala 475:29]
  reg  bus_cmd_req_hold; // @[Reg.scala 27:20]
  wire  _T_2617 = ic_act_miss_f | bus_cmd_req_hold; // @[ifu_mem_ctl.scala 462:45]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2618 = _T_2617 | ifu_bus_cmd_valid; // @[ifu_mem_ctl.scala 462:64]
  wire  _T_2620 = _T_2618 & _T_2653; // @[ifu_mem_ctl.scala 462:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2622 = bus_cmd_beat_count == 3'h7; // @[ifu_mem_ctl.scala 462:146]
  wire  _T_2623 = _T_2622 & ifu_bus_cmd_valid; // @[ifu_mem_ctl.scala 462:177]
  wire  _T_2624 = _T_2623 & io_ifu_axi_ar_ready; // @[ifu_mem_ctl.scala 462:197]
  wire  _T_2625 = _T_2624 & miss_pending; // @[ifu_mem_ctl.scala 462:219]
  wire  _T_2626 = ~_T_2625; // @[ifu_mem_ctl.scala 462:125]
  wire  ifc_bus_ic_req_ff_in = _T_2620 & _T_2626; // @[ifu_mem_ctl.scala 462:123]
  wire  _T_2627 = io_ifu_bus_clk_en | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 463:88]
  wire  ifu_bus_arready = io_ifu_axi_ar_ready & io_ifu_bus_clk_en; // @[ifu_mem_ctl.scala 486:45]
  wire  _T_2647 = io_ifu_axi_ar_valid & ifu_bus_arready; // @[ifu_mem_ctl.scala 490:39]
  wire  _T_2648 = _T_2647 & miss_pending; // @[ifu_mem_ctl.scala 490:57]
  wire  bus_cmd_sent = _T_2648 & _T_2653; // @[ifu_mem_ctl.scala 490:72]
  wire  _T_2630 = ~bus_cmd_sent; // @[ifu_mem_ctl.scala 465:61]
  wire  _T_2631 = _T_2617 & _T_2630; // @[ifu_mem_ctl.scala 465:59]
  wire  bus_cmd_req_in = _T_2631 & _T_2653; // @[ifu_mem_ctl.scala 465:75]
  wire  _T_2634 = bus_cmd_req_in ^ bus_cmd_req_hold; // @[lib.scala 475:21]
  wire  _T_2635 = |_T_2634; // @[lib.scala 475:29]
  wire [2:0] _T_2639 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2641 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2643 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[ifu_mem_ctl.scala 487:51]
  wire [2:0] _T_2667 = bus_new_data_beat_count ^ bus_data_beat_count; // @[lib.scala 453:21]
  wire  _T_2668 = |_T_2667; // @[lib.scala 453:29]
  wire  _T_2671 = ~scnd_miss_req; // @[ifu_mem_ctl.scala 498:73]
  wire  _T_2672 = _T_2654 & _T_2671; // @[ifu_mem_ctl.scala 498:71]
  wire  _T_2674 = last_data_recieved_ff & _T_1362; // @[ifu_mem_ctl.scala 498:114]
  wire  last_data_recieved_in = _T_2672 | _T_2674; // @[ifu_mem_ctl.scala 498:89]
  wire  _T_2676 = last_data_recieved_in ^ last_data_recieved_ff; // @[lib.scala 475:21]
  wire  _T_2677 = |_T_2676; // @[lib.scala 475:29]
  wire [2:0] _T_2683 = bus_rd_addr_count + 3'h1; // @[ifu_mem_ctl.scala 503:43]
  wire  _T_2689 = ifu_bus_cmd_valid & io_ifu_axi_ar_ready; // @[ifu_mem_ctl.scala 506:48]
  wire  _T_2690 = _T_2689 & miss_pending; // @[ifu_mem_ctl.scala 506:70]
  wire  bus_inc_cmd_beat_cnt = _T_2690 & _T_2653; // @[ifu_mem_ctl.scala 506:85]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[ifu_mem_ctl.scala 508:57]
  wire  _T_2694 = ~bus_inc_cmd_beat_cnt; // @[ifu_mem_ctl.scala 509:31]
  wire  _T_2695 = ic_act_miss_f | scnd_miss_req; // @[ifu_mem_ctl.scala 509:71]
  wire  _T_2696 = _T_2695 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 509:87]
  wire  _T_2697 = ~_T_2696; // @[ifu_mem_ctl.scala 509:55]
  wire  bus_hold_cmd_beat_cnt = _T_2694 & _T_2697; // @[ifu_mem_ctl.scala 509:53]
  wire  _T_2698 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[ifu_mem_ctl.scala 510:46]
  wire  bus_cmd_beat_en = _T_2698 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 510:62]
  wire [2:0] _T_2701 = bus_cmd_beat_count + 3'h1; // @[ifu_mem_ctl.scala 512:46]
  wire [2:0] _T_2703 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2704 = bus_inc_cmd_beat_cnt ? _T_2701 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2705 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2707 = _T_2703 | _T_2704; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2707 | _T_2705; // @[Mux.scala 27:72]
  wire  _T_2711 = _T_326 & bus_cmd_beat_en; // @[lib.scala 393:57]
  wire  _T_2727 = ic_act_miss_f ^ ic_act_miss_f_delayed; // @[lib.scala 475:21]
  wire  _T_2728 = |_T_2727; // @[lib.scala 475:29]
  wire  _T_2740 = ~iccm_correct_ecc; // @[ifu_mem_ctl.scala 523:53]
  wire  _T_2741 = io_ifc_dma_access_ok & _T_2740; // @[ifu_mem_ctl.scala 523:50]
  wire  _T_2742 = ~io_iccm_dma_sb_error; // @[ifu_mem_ctl.scala 523:73]
  wire  ifc_dma_access_ok_d = _T_2741 & _T_2742; // @[ifu_mem_ctl.scala 523:71]
  reg  ifc_dma_access_ok_prev; // @[Reg.scala 27:20]
  wire  _T_2743 = ifc_dma_access_ok_d ^ ifc_dma_access_ok_prev; // @[lib.scala 475:21]
  wire  _T_2744 = |_T_2743; // @[lib.scala 475:29]
  wire  _T_2750 = _T_2741 & ifc_dma_access_ok_prev; // @[ifu_mem_ctl.scala 530:63]
  wire  _T_2751 = perr_state == 3'h0; // @[ifu_mem_ctl.scala 530:102]
  wire  _T_2752 = _T_2750 & _T_2751; // @[ifu_mem_ctl.scala 530:88]
  wire  _T_2756 = io_dma_mem_ctl_dma_iccm_req ^ dma_iccm_req_f; // @[lib.scala 475:21]
  wire  _T_2757 = |_T_2756; // @[lib.scala 475:29]
  wire  _T_2759 = io_iccm_ready & io_dma_mem_ctl_dma_iccm_req; // @[ifu_mem_ctl.scala 532:34]
  wire  _T_2760 = _T_2759 & io_dma_mem_ctl_dma_mem_write; // @[ifu_mem_ctl.scala 532:64]
  wire  _T_2763 = ~io_dma_mem_ctl_dma_mem_write; // @[ifu_mem_ctl.scala 533:66]
  wire  _T_2764 = _T_2759 & _T_2763; // @[ifu_mem_ctl.scala 533:64]
  wire  _T_2765 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[ifu_mem_ctl.scala 533:122]
  wire [2:0] _T_2770 = io_dma_mem_ctl_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire  _T_2791 = io_dma_mem_ctl_dma_mem_wdata[32] ^ io_dma_mem_ctl_dma_mem_wdata[33]; // @[lib.scala 119:74]
  wire  _T_2792 = _T_2791 ^ io_dma_mem_ctl_dma_mem_wdata[35]; // @[lib.scala 119:74]
  wire  _T_2793 = _T_2792 ^ io_dma_mem_ctl_dma_mem_wdata[36]; // @[lib.scala 119:74]
  wire  _T_2794 = _T_2793 ^ io_dma_mem_ctl_dma_mem_wdata[38]; // @[lib.scala 119:74]
  wire  _T_2795 = _T_2794 ^ io_dma_mem_ctl_dma_mem_wdata[40]; // @[lib.scala 119:74]
  wire  _T_2796 = _T_2795 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2797 = _T_2796 ^ io_dma_mem_ctl_dma_mem_wdata[43]; // @[lib.scala 119:74]
  wire  _T_2798 = _T_2797 ^ io_dma_mem_ctl_dma_mem_wdata[45]; // @[lib.scala 119:74]
  wire  _T_2799 = _T_2798 ^ io_dma_mem_ctl_dma_mem_wdata[47]; // @[lib.scala 119:74]
  wire  _T_2800 = _T_2799 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2801 = _T_2800 ^ io_dma_mem_ctl_dma_mem_wdata[51]; // @[lib.scala 119:74]
  wire  _T_2802 = _T_2801 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2803 = _T_2802 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2804 = _T_2803 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2805 = _T_2804 ^ io_dma_mem_ctl_dma_mem_wdata[58]; // @[lib.scala 119:74]
  wire  _T_2806 = _T_2805 ^ io_dma_mem_ctl_dma_mem_wdata[60]; // @[lib.scala 119:74]
  wire  _T_2807 = _T_2806 ^ io_dma_mem_ctl_dma_mem_wdata[62]; // @[lib.scala 119:74]
  wire  _T_2826 = io_dma_mem_ctl_dma_mem_wdata[32] ^ io_dma_mem_ctl_dma_mem_wdata[34]; // @[lib.scala 119:74]
  wire  _T_2827 = _T_2826 ^ io_dma_mem_ctl_dma_mem_wdata[35]; // @[lib.scala 119:74]
  wire  _T_2828 = _T_2827 ^ io_dma_mem_ctl_dma_mem_wdata[37]; // @[lib.scala 119:74]
  wire  _T_2829 = _T_2828 ^ io_dma_mem_ctl_dma_mem_wdata[38]; // @[lib.scala 119:74]
  wire  _T_2830 = _T_2829 ^ io_dma_mem_ctl_dma_mem_wdata[41]; // @[lib.scala 119:74]
  wire  _T_2831 = _T_2830 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2832 = _T_2831 ^ io_dma_mem_ctl_dma_mem_wdata[44]; // @[lib.scala 119:74]
  wire  _T_2833 = _T_2832 ^ io_dma_mem_ctl_dma_mem_wdata[45]; // @[lib.scala 119:74]
  wire  _T_2834 = _T_2833 ^ io_dma_mem_ctl_dma_mem_wdata[48]; // @[lib.scala 119:74]
  wire  _T_2835 = _T_2834 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2836 = _T_2835 ^ io_dma_mem_ctl_dma_mem_wdata[52]; // @[lib.scala 119:74]
  wire  _T_2837 = _T_2836 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2838 = _T_2837 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2839 = _T_2838 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2840 = _T_2839 ^ io_dma_mem_ctl_dma_mem_wdata[59]; // @[lib.scala 119:74]
  wire  _T_2841 = _T_2840 ^ io_dma_mem_ctl_dma_mem_wdata[60]; // @[lib.scala 119:74]
  wire  _T_2842 = _T_2841 ^ io_dma_mem_ctl_dma_mem_wdata[63]; // @[lib.scala 119:74]
  wire  _T_2861 = io_dma_mem_ctl_dma_mem_wdata[33] ^ io_dma_mem_ctl_dma_mem_wdata[34]; // @[lib.scala 119:74]
  wire  _T_2862 = _T_2861 ^ io_dma_mem_ctl_dma_mem_wdata[35]; // @[lib.scala 119:74]
  wire  _T_2863 = _T_2862 ^ io_dma_mem_ctl_dma_mem_wdata[39]; // @[lib.scala 119:74]
  wire  _T_2864 = _T_2863 ^ io_dma_mem_ctl_dma_mem_wdata[40]; // @[lib.scala 119:74]
  wire  _T_2865 = _T_2864 ^ io_dma_mem_ctl_dma_mem_wdata[41]; // @[lib.scala 119:74]
  wire  _T_2866 = _T_2865 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2867 = _T_2866 ^ io_dma_mem_ctl_dma_mem_wdata[46]; // @[lib.scala 119:74]
  wire  _T_2868 = _T_2867 ^ io_dma_mem_ctl_dma_mem_wdata[47]; // @[lib.scala 119:74]
  wire  _T_2869 = _T_2868 ^ io_dma_mem_ctl_dma_mem_wdata[48]; // @[lib.scala 119:74]
  wire  _T_2870 = _T_2869 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2871 = _T_2870 ^ io_dma_mem_ctl_dma_mem_wdata[54]; // @[lib.scala 119:74]
  wire  _T_2872 = _T_2871 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2873 = _T_2872 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2874 = _T_2873 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2875 = _T_2874 ^ io_dma_mem_ctl_dma_mem_wdata[61]; // @[lib.scala 119:74]
  wire  _T_2876 = _T_2875 ^ io_dma_mem_ctl_dma_mem_wdata[62]; // @[lib.scala 119:74]
  wire  _T_2877 = _T_2876 ^ io_dma_mem_ctl_dma_mem_wdata[63]; // @[lib.scala 119:74]
  wire  _T_2893 = io_dma_mem_ctl_dma_mem_wdata[36] ^ io_dma_mem_ctl_dma_mem_wdata[37]; // @[lib.scala 119:74]
  wire  _T_2894 = _T_2893 ^ io_dma_mem_ctl_dma_mem_wdata[38]; // @[lib.scala 119:74]
  wire  _T_2895 = _T_2894 ^ io_dma_mem_ctl_dma_mem_wdata[39]; // @[lib.scala 119:74]
  wire  _T_2896 = _T_2895 ^ io_dma_mem_ctl_dma_mem_wdata[40]; // @[lib.scala 119:74]
  wire  _T_2897 = _T_2896 ^ io_dma_mem_ctl_dma_mem_wdata[41]; // @[lib.scala 119:74]
  wire  _T_2898 = _T_2897 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2899 = _T_2898 ^ io_dma_mem_ctl_dma_mem_wdata[50]; // @[lib.scala 119:74]
  wire  _T_2900 = _T_2899 ^ io_dma_mem_ctl_dma_mem_wdata[51]; // @[lib.scala 119:74]
  wire  _T_2901 = _T_2900 ^ io_dma_mem_ctl_dma_mem_wdata[52]; // @[lib.scala 119:74]
  wire  _T_2902 = _T_2901 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2903 = _T_2902 ^ io_dma_mem_ctl_dma_mem_wdata[54]; // @[lib.scala 119:74]
  wire  _T_2904 = _T_2903 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2905 = _T_2904 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2906 = _T_2905 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2922 = io_dma_mem_ctl_dma_mem_wdata[43] ^ io_dma_mem_ctl_dma_mem_wdata[44]; // @[lib.scala 119:74]
  wire  _T_2923 = _T_2922 ^ io_dma_mem_ctl_dma_mem_wdata[45]; // @[lib.scala 119:74]
  wire  _T_2924 = _T_2923 ^ io_dma_mem_ctl_dma_mem_wdata[46]; // @[lib.scala 119:74]
  wire  _T_2925 = _T_2924 ^ io_dma_mem_ctl_dma_mem_wdata[47]; // @[lib.scala 119:74]
  wire  _T_2926 = _T_2925 ^ io_dma_mem_ctl_dma_mem_wdata[48]; // @[lib.scala 119:74]
  wire  _T_2927 = _T_2926 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2928 = _T_2927 ^ io_dma_mem_ctl_dma_mem_wdata[50]; // @[lib.scala 119:74]
  wire  _T_2929 = _T_2928 ^ io_dma_mem_ctl_dma_mem_wdata[51]; // @[lib.scala 119:74]
  wire  _T_2930 = _T_2929 ^ io_dma_mem_ctl_dma_mem_wdata[52]; // @[lib.scala 119:74]
  wire  _T_2931 = _T_2930 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2932 = _T_2931 ^ io_dma_mem_ctl_dma_mem_wdata[54]; // @[lib.scala 119:74]
  wire  _T_2933 = _T_2932 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2934 = _T_2933 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2935 = _T_2934 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2942 = io_dma_mem_ctl_dma_mem_wdata[58] ^ io_dma_mem_ctl_dma_mem_wdata[59]; // @[lib.scala 119:74]
  wire  _T_2943 = _T_2942 ^ io_dma_mem_ctl_dma_mem_wdata[60]; // @[lib.scala 119:74]
  wire  _T_2944 = _T_2943 ^ io_dma_mem_ctl_dma_mem_wdata[61]; // @[lib.scala 119:74]
  wire  _T_2945 = _T_2944 ^ io_dma_mem_ctl_dma_mem_wdata[62]; // @[lib.scala 119:74]
  wire  _T_2946 = _T_2945 ^ io_dma_mem_ctl_dma_mem_wdata[63]; // @[lib.scala 119:74]
  wire [5:0] _T_2951 = {_T_2946,_T_2935,_T_2906,_T_2877,_T_2842,_T_2807}; // @[Cat.scala 29:58]
  wire  _T_2952 = ^io_dma_mem_ctl_dma_mem_wdata[63:32]; // @[lib.scala 127:13]
  wire  _T_2953 = ^_T_2951; // @[lib.scala 127:23]
  wire  _T_2954 = _T_2952 ^ _T_2953; // @[lib.scala 127:18]
  wire  _T_2975 = io_dma_mem_ctl_dma_mem_wdata[0] ^ io_dma_mem_ctl_dma_mem_wdata[1]; // @[lib.scala 119:74]
  wire  _T_2976 = _T_2975 ^ io_dma_mem_ctl_dma_mem_wdata[3]; // @[lib.scala 119:74]
  wire  _T_2977 = _T_2976 ^ io_dma_mem_ctl_dma_mem_wdata[4]; // @[lib.scala 119:74]
  wire  _T_2978 = _T_2977 ^ io_dma_mem_ctl_dma_mem_wdata[6]; // @[lib.scala 119:74]
  wire  _T_2979 = _T_2978 ^ io_dma_mem_ctl_dma_mem_wdata[8]; // @[lib.scala 119:74]
  wire  _T_2980 = _T_2979 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_2981 = _T_2980 ^ io_dma_mem_ctl_dma_mem_wdata[11]; // @[lib.scala 119:74]
  wire  _T_2982 = _T_2981 ^ io_dma_mem_ctl_dma_mem_wdata[13]; // @[lib.scala 119:74]
  wire  _T_2983 = _T_2982 ^ io_dma_mem_ctl_dma_mem_wdata[15]; // @[lib.scala 119:74]
  wire  _T_2984 = _T_2983 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_2985 = _T_2984 ^ io_dma_mem_ctl_dma_mem_wdata[19]; // @[lib.scala 119:74]
  wire  _T_2986 = _T_2985 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_2987 = _T_2986 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_2988 = _T_2987 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_2989 = _T_2988 ^ io_dma_mem_ctl_dma_mem_wdata[26]; // @[lib.scala 119:74]
  wire  _T_2990 = _T_2989 ^ io_dma_mem_ctl_dma_mem_wdata[28]; // @[lib.scala 119:74]
  wire  _T_2991 = _T_2990 ^ io_dma_mem_ctl_dma_mem_wdata[30]; // @[lib.scala 119:74]
  wire  _T_3010 = io_dma_mem_ctl_dma_mem_wdata[0] ^ io_dma_mem_ctl_dma_mem_wdata[2]; // @[lib.scala 119:74]
  wire  _T_3011 = _T_3010 ^ io_dma_mem_ctl_dma_mem_wdata[3]; // @[lib.scala 119:74]
  wire  _T_3012 = _T_3011 ^ io_dma_mem_ctl_dma_mem_wdata[5]; // @[lib.scala 119:74]
  wire  _T_3013 = _T_3012 ^ io_dma_mem_ctl_dma_mem_wdata[6]; // @[lib.scala 119:74]
  wire  _T_3014 = _T_3013 ^ io_dma_mem_ctl_dma_mem_wdata[9]; // @[lib.scala 119:74]
  wire  _T_3015 = _T_3014 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_3016 = _T_3015 ^ io_dma_mem_ctl_dma_mem_wdata[12]; // @[lib.scala 119:74]
  wire  _T_3017 = _T_3016 ^ io_dma_mem_ctl_dma_mem_wdata[13]; // @[lib.scala 119:74]
  wire  _T_3018 = _T_3017 ^ io_dma_mem_ctl_dma_mem_wdata[16]; // @[lib.scala 119:74]
  wire  _T_3019 = _T_3018 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_3020 = _T_3019 ^ io_dma_mem_ctl_dma_mem_wdata[20]; // @[lib.scala 119:74]
  wire  _T_3021 = _T_3020 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_3022 = _T_3021 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_3023 = _T_3022 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_3024 = _T_3023 ^ io_dma_mem_ctl_dma_mem_wdata[27]; // @[lib.scala 119:74]
  wire  _T_3025 = _T_3024 ^ io_dma_mem_ctl_dma_mem_wdata[28]; // @[lib.scala 119:74]
  wire  _T_3026 = _T_3025 ^ io_dma_mem_ctl_dma_mem_wdata[31]; // @[lib.scala 119:74]
  wire  _T_3045 = io_dma_mem_ctl_dma_mem_wdata[1] ^ io_dma_mem_ctl_dma_mem_wdata[2]; // @[lib.scala 119:74]
  wire  _T_3046 = _T_3045 ^ io_dma_mem_ctl_dma_mem_wdata[3]; // @[lib.scala 119:74]
  wire  _T_3047 = _T_3046 ^ io_dma_mem_ctl_dma_mem_wdata[7]; // @[lib.scala 119:74]
  wire  _T_3048 = _T_3047 ^ io_dma_mem_ctl_dma_mem_wdata[8]; // @[lib.scala 119:74]
  wire  _T_3049 = _T_3048 ^ io_dma_mem_ctl_dma_mem_wdata[9]; // @[lib.scala 119:74]
  wire  _T_3050 = _T_3049 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_3051 = _T_3050 ^ io_dma_mem_ctl_dma_mem_wdata[14]; // @[lib.scala 119:74]
  wire  _T_3052 = _T_3051 ^ io_dma_mem_ctl_dma_mem_wdata[15]; // @[lib.scala 119:74]
  wire  _T_3053 = _T_3052 ^ io_dma_mem_ctl_dma_mem_wdata[16]; // @[lib.scala 119:74]
  wire  _T_3054 = _T_3053 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_3055 = _T_3054 ^ io_dma_mem_ctl_dma_mem_wdata[22]; // @[lib.scala 119:74]
  wire  _T_3056 = _T_3055 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_3057 = _T_3056 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_3058 = _T_3057 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_3059 = _T_3058 ^ io_dma_mem_ctl_dma_mem_wdata[29]; // @[lib.scala 119:74]
  wire  _T_3060 = _T_3059 ^ io_dma_mem_ctl_dma_mem_wdata[30]; // @[lib.scala 119:74]
  wire  _T_3061 = _T_3060 ^ io_dma_mem_ctl_dma_mem_wdata[31]; // @[lib.scala 119:74]
  wire  _T_3077 = io_dma_mem_ctl_dma_mem_wdata[4] ^ io_dma_mem_ctl_dma_mem_wdata[5]; // @[lib.scala 119:74]
  wire  _T_3078 = _T_3077 ^ io_dma_mem_ctl_dma_mem_wdata[6]; // @[lib.scala 119:74]
  wire  _T_3079 = _T_3078 ^ io_dma_mem_ctl_dma_mem_wdata[7]; // @[lib.scala 119:74]
  wire  _T_3080 = _T_3079 ^ io_dma_mem_ctl_dma_mem_wdata[8]; // @[lib.scala 119:74]
  wire  _T_3081 = _T_3080 ^ io_dma_mem_ctl_dma_mem_wdata[9]; // @[lib.scala 119:74]
  wire  _T_3082 = _T_3081 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_3083 = _T_3082 ^ io_dma_mem_ctl_dma_mem_wdata[18]; // @[lib.scala 119:74]
  wire  _T_3084 = _T_3083 ^ io_dma_mem_ctl_dma_mem_wdata[19]; // @[lib.scala 119:74]
  wire  _T_3085 = _T_3084 ^ io_dma_mem_ctl_dma_mem_wdata[20]; // @[lib.scala 119:74]
  wire  _T_3086 = _T_3085 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_3087 = _T_3086 ^ io_dma_mem_ctl_dma_mem_wdata[22]; // @[lib.scala 119:74]
  wire  _T_3088 = _T_3087 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_3089 = _T_3088 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_3090 = _T_3089 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_3106 = io_dma_mem_ctl_dma_mem_wdata[11] ^ io_dma_mem_ctl_dma_mem_wdata[12]; // @[lib.scala 119:74]
  wire  _T_3107 = _T_3106 ^ io_dma_mem_ctl_dma_mem_wdata[13]; // @[lib.scala 119:74]
  wire  _T_3108 = _T_3107 ^ io_dma_mem_ctl_dma_mem_wdata[14]; // @[lib.scala 119:74]
  wire  _T_3109 = _T_3108 ^ io_dma_mem_ctl_dma_mem_wdata[15]; // @[lib.scala 119:74]
  wire  _T_3110 = _T_3109 ^ io_dma_mem_ctl_dma_mem_wdata[16]; // @[lib.scala 119:74]
  wire  _T_3111 = _T_3110 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_3112 = _T_3111 ^ io_dma_mem_ctl_dma_mem_wdata[18]; // @[lib.scala 119:74]
  wire  _T_3113 = _T_3112 ^ io_dma_mem_ctl_dma_mem_wdata[19]; // @[lib.scala 119:74]
  wire  _T_3114 = _T_3113 ^ io_dma_mem_ctl_dma_mem_wdata[20]; // @[lib.scala 119:74]
  wire  _T_3115 = _T_3114 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_3116 = _T_3115 ^ io_dma_mem_ctl_dma_mem_wdata[22]; // @[lib.scala 119:74]
  wire  _T_3117 = _T_3116 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_3118 = _T_3117 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_3119 = _T_3118 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_3126 = io_dma_mem_ctl_dma_mem_wdata[26] ^ io_dma_mem_ctl_dma_mem_wdata[27]; // @[lib.scala 119:74]
  wire  _T_3127 = _T_3126 ^ io_dma_mem_ctl_dma_mem_wdata[28]; // @[lib.scala 119:74]
  wire  _T_3128 = _T_3127 ^ io_dma_mem_ctl_dma_mem_wdata[29]; // @[lib.scala 119:74]
  wire  _T_3129 = _T_3128 ^ io_dma_mem_ctl_dma_mem_wdata[30]; // @[lib.scala 119:74]
  wire  _T_3130 = _T_3129 ^ io_dma_mem_ctl_dma_mem_wdata[31]; // @[lib.scala 119:74]
  wire [5:0] _T_3135 = {_T_3130,_T_3119,_T_3090,_T_3061,_T_3026,_T_2991}; // @[Cat.scala 29:58]
  wire  _T_3136 = ^io_dma_mem_ctl_dma_mem_wdata[31:0]; // @[lib.scala 127:13]
  wire  _T_3137 = ^_T_3135; // @[lib.scala 127:23]
  wire  _T_3138 = _T_3136 ^ _T_3137; // @[lib.scala 127:18]
  wire [6:0] _T_3139 = {_T_3138,_T_3130,_T_3119,_T_3090,_T_3061,_T_3026,_T_2991}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2954,_T_2946,_T_2935,_T_2906,_T_2877,_T_2842,_T_2807,_T_3139}; // @[Cat.scala 29:58]
  wire  _T_3141 = ~_T_2759; // @[ifu_mem_ctl.scala 539:45]
  wire  _T_3142 = iccm_correct_ecc & _T_3141; // @[ifu_mem_ctl.scala 539:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3143 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3150 = {dma_mem_ecc[13:7],io_dma_mem_ctl_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_ctl_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[Reg.scala 27:20]
  wire  _T_3505 = _T_3417[5:0] == 6'h27; // @[lib.scala 199:41]
  wire  _T_3503 = _T_3417[5:0] == 6'h26; // @[lib.scala 199:41]
  wire  _T_3501 = _T_3417[5:0] == 6'h25; // @[lib.scala 199:41]
  wire  _T_3499 = _T_3417[5:0] == 6'h24; // @[lib.scala 199:41]
  wire  _T_3497 = _T_3417[5:0] == 6'h23; // @[lib.scala 199:41]
  wire  _T_3495 = _T_3417[5:0] == 6'h22; // @[lib.scala 199:41]
  wire  _T_3493 = _T_3417[5:0] == 6'h21; // @[lib.scala 199:41]
  wire  _T_3491 = _T_3417[5:0] == 6'h20; // @[lib.scala 199:41]
  wire  _T_3489 = _T_3417[5:0] == 6'h1f; // @[lib.scala 199:41]
  wire  _T_3487 = _T_3417[5:0] == 6'h1e; // @[lib.scala 199:41]
  wire [9:0] _T_3563 = {_T_3505,_T_3503,_T_3501,_T_3499,_T_3497,_T_3495,_T_3493,_T_3491,_T_3489,_T_3487}; // @[lib.scala 202:69]
  wire  _T_3485 = _T_3417[5:0] == 6'h1d; // @[lib.scala 199:41]
  wire  _T_3483 = _T_3417[5:0] == 6'h1c; // @[lib.scala 199:41]
  wire  _T_3481 = _T_3417[5:0] == 6'h1b; // @[lib.scala 199:41]
  wire  _T_3479 = _T_3417[5:0] == 6'h1a; // @[lib.scala 199:41]
  wire  _T_3477 = _T_3417[5:0] == 6'h19; // @[lib.scala 199:41]
  wire  _T_3475 = _T_3417[5:0] == 6'h18; // @[lib.scala 199:41]
  wire  _T_3473 = _T_3417[5:0] == 6'h17; // @[lib.scala 199:41]
  wire  _T_3471 = _T_3417[5:0] == 6'h16; // @[lib.scala 199:41]
  wire  _T_3469 = _T_3417[5:0] == 6'h15; // @[lib.scala 199:41]
  wire  _T_3467 = _T_3417[5:0] == 6'h14; // @[lib.scala 199:41]
  wire [9:0] _T_3554 = {_T_3485,_T_3483,_T_3481,_T_3479,_T_3477,_T_3475,_T_3473,_T_3471,_T_3469,_T_3467}; // @[lib.scala 202:69]
  wire  _T_3465 = _T_3417[5:0] == 6'h13; // @[lib.scala 199:41]
  wire  _T_3463 = _T_3417[5:0] == 6'h12; // @[lib.scala 199:41]
  wire  _T_3461 = _T_3417[5:0] == 6'h11; // @[lib.scala 199:41]
  wire  _T_3459 = _T_3417[5:0] == 6'h10; // @[lib.scala 199:41]
  wire  _T_3457 = _T_3417[5:0] == 6'hf; // @[lib.scala 199:41]
  wire  _T_3455 = _T_3417[5:0] == 6'he; // @[lib.scala 199:41]
  wire  _T_3453 = _T_3417[5:0] == 6'hd; // @[lib.scala 199:41]
  wire  _T_3451 = _T_3417[5:0] == 6'hc; // @[lib.scala 199:41]
  wire  _T_3449 = _T_3417[5:0] == 6'hb; // @[lib.scala 199:41]
  wire  _T_3447 = _T_3417[5:0] == 6'ha; // @[lib.scala 199:41]
  wire [9:0] _T_3544 = {_T_3465,_T_3463,_T_3461,_T_3459,_T_3457,_T_3455,_T_3453,_T_3451,_T_3449,_T_3447}; // @[lib.scala 202:69]
  wire  _T_3445 = _T_3417[5:0] == 6'h9; // @[lib.scala 199:41]
  wire  _T_3443 = _T_3417[5:0] == 6'h8; // @[lib.scala 199:41]
  wire  _T_3441 = _T_3417[5:0] == 6'h7; // @[lib.scala 199:41]
  wire  _T_3439 = _T_3417[5:0] == 6'h6; // @[lib.scala 199:41]
  wire  _T_3437 = _T_3417[5:0] == 6'h5; // @[lib.scala 199:41]
  wire  _T_3435 = _T_3417[5:0] == 6'h4; // @[lib.scala 199:41]
  wire  _T_3433 = _T_3417[5:0] == 6'h3; // @[lib.scala 199:41]
  wire  _T_3431 = _T_3417[5:0] == 6'h2; // @[lib.scala 199:41]
  wire  _T_3429 = _T_3417[5:0] == 6'h1; // @[lib.scala 199:41]
  wire [18:0] _T_3545 = {_T_3544,_T_3445,_T_3443,_T_3441,_T_3439,_T_3437,_T_3435,_T_3433,_T_3431,_T_3429}; // @[lib.scala 202:69]
  wire [38:0] _T_3565 = {_T_3563,_T_3554,_T_3545}; // @[lib.scala 202:69]
  wire [7:0] _T_3520 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3526 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3520}; // @[Cat.scala 29:58]
  wire [38:0] _T_3566 = _T_3565 ^ _T_3526; // @[lib.scala 202:76]
  wire [38:0] _T_3567 = _T_3421 ? _T_3566 : _T_3526; // @[lib.scala 202:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3567[37:32],_T_3567[30:16],_T_3567[14:8],_T_3567[6:4],_T_3567[2]}; // @[Cat.scala 29:58]
  wire  _T_3890 = _T_3802[5:0] == 6'h27; // @[lib.scala 199:41]
  wire  _T_3888 = _T_3802[5:0] == 6'h26; // @[lib.scala 199:41]
  wire  _T_3886 = _T_3802[5:0] == 6'h25; // @[lib.scala 199:41]
  wire  _T_3884 = _T_3802[5:0] == 6'h24; // @[lib.scala 199:41]
  wire  _T_3882 = _T_3802[5:0] == 6'h23; // @[lib.scala 199:41]
  wire  _T_3880 = _T_3802[5:0] == 6'h22; // @[lib.scala 199:41]
  wire  _T_3878 = _T_3802[5:0] == 6'h21; // @[lib.scala 199:41]
  wire  _T_3876 = _T_3802[5:0] == 6'h20; // @[lib.scala 199:41]
  wire  _T_3874 = _T_3802[5:0] == 6'h1f; // @[lib.scala 199:41]
  wire  _T_3872 = _T_3802[5:0] == 6'h1e; // @[lib.scala 199:41]
  wire [9:0] _T_3948 = {_T_3890,_T_3888,_T_3886,_T_3884,_T_3882,_T_3880,_T_3878,_T_3876,_T_3874,_T_3872}; // @[lib.scala 202:69]
  wire  _T_3870 = _T_3802[5:0] == 6'h1d; // @[lib.scala 199:41]
  wire  _T_3868 = _T_3802[5:0] == 6'h1c; // @[lib.scala 199:41]
  wire  _T_3866 = _T_3802[5:0] == 6'h1b; // @[lib.scala 199:41]
  wire  _T_3864 = _T_3802[5:0] == 6'h1a; // @[lib.scala 199:41]
  wire  _T_3862 = _T_3802[5:0] == 6'h19; // @[lib.scala 199:41]
  wire  _T_3860 = _T_3802[5:0] == 6'h18; // @[lib.scala 199:41]
  wire  _T_3858 = _T_3802[5:0] == 6'h17; // @[lib.scala 199:41]
  wire  _T_3856 = _T_3802[5:0] == 6'h16; // @[lib.scala 199:41]
  wire  _T_3854 = _T_3802[5:0] == 6'h15; // @[lib.scala 199:41]
  wire  _T_3852 = _T_3802[5:0] == 6'h14; // @[lib.scala 199:41]
  wire [9:0] _T_3939 = {_T_3870,_T_3868,_T_3866,_T_3864,_T_3862,_T_3860,_T_3858,_T_3856,_T_3854,_T_3852}; // @[lib.scala 202:69]
  wire  _T_3850 = _T_3802[5:0] == 6'h13; // @[lib.scala 199:41]
  wire  _T_3848 = _T_3802[5:0] == 6'h12; // @[lib.scala 199:41]
  wire  _T_3846 = _T_3802[5:0] == 6'h11; // @[lib.scala 199:41]
  wire  _T_3844 = _T_3802[5:0] == 6'h10; // @[lib.scala 199:41]
  wire  _T_3842 = _T_3802[5:0] == 6'hf; // @[lib.scala 199:41]
  wire  _T_3840 = _T_3802[5:0] == 6'he; // @[lib.scala 199:41]
  wire  _T_3838 = _T_3802[5:0] == 6'hd; // @[lib.scala 199:41]
  wire  _T_3836 = _T_3802[5:0] == 6'hc; // @[lib.scala 199:41]
  wire  _T_3834 = _T_3802[5:0] == 6'hb; // @[lib.scala 199:41]
  wire  _T_3832 = _T_3802[5:0] == 6'ha; // @[lib.scala 199:41]
  wire [9:0] _T_3929 = {_T_3850,_T_3848,_T_3846,_T_3844,_T_3842,_T_3840,_T_3838,_T_3836,_T_3834,_T_3832}; // @[lib.scala 202:69]
  wire  _T_3830 = _T_3802[5:0] == 6'h9; // @[lib.scala 199:41]
  wire  _T_3828 = _T_3802[5:0] == 6'h8; // @[lib.scala 199:41]
  wire  _T_3826 = _T_3802[5:0] == 6'h7; // @[lib.scala 199:41]
  wire  _T_3824 = _T_3802[5:0] == 6'h6; // @[lib.scala 199:41]
  wire  _T_3822 = _T_3802[5:0] == 6'h5; // @[lib.scala 199:41]
  wire  _T_3820 = _T_3802[5:0] == 6'h4; // @[lib.scala 199:41]
  wire  _T_3818 = _T_3802[5:0] == 6'h3; // @[lib.scala 199:41]
  wire  _T_3816 = _T_3802[5:0] == 6'h2; // @[lib.scala 199:41]
  wire  _T_3814 = _T_3802[5:0] == 6'h1; // @[lib.scala 199:41]
  wire [18:0] _T_3930 = {_T_3929,_T_3830,_T_3828,_T_3826,_T_3824,_T_3822,_T_3820,_T_3818,_T_3816,_T_3814}; // @[lib.scala 202:69]
  wire [38:0] _T_3950 = {_T_3948,_T_3939,_T_3930}; // @[lib.scala 202:69]
  wire [7:0] _T_3905 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3911 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3905}; // @[Cat.scala 29:58]
  wire [38:0] _T_3951 = _T_3950 ^ _T_3911; // @[lib.scala 202:76]
  wire [38:0] _T_3952 = _T_3806 ? _T_3951 : _T_3911; // @[lib.scala 202:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3952[37:32],_T_3952[30:16],_T_3952[14:8],_T_3952[6:4],_T_3952[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[ifu_mem_ctl.scala 543:35]
  wire  _T_3810 = ~_T_3802[6]; // @[lib.scala 195:55]
  wire  _T_3811 = _T_3804 & _T_3810; // @[lib.scala 195:53]
  wire  _T_3425 = ~_T_3417[6]; // @[lib.scala 195:55]
  wire  _T_3426 = _T_3419 & _T_3425; // @[lib.scala 195:53]
  wire [1:0] iccm_double_ecc_error = {_T_3811,_T_3426}; // @[Cat.scala 29:58]
  wire  _T_3154 = |iccm_double_ecc_error; // @[ifu_mem_ctl.scala 545:53]
  wire [63:0] _T_3155 = {io_dma_mem_ctl_dma_mem_addr,io_dma_mem_ctl_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3156 = {iccm_dma_rdata_1_muxed,_T_3567[37:32],_T_3567[30:16],_T_3567[14:8],_T_3567[6:4],_T_3567[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[Reg.scala 27:20]
  wire [2:0] _T_3157 = io_dma_mem_ctl_dma_mem_tag ^ dma_mem_tag_ff; // @[lib.scala 453:21]
  wire  _T_3158 = |_T_3157; // @[lib.scala 453:29]
  reg [2:0] iccm_dma_rtag_temp; // @[Reg.scala 27:20]
  wire [2:0] _T_3160 = dma_mem_tag_ff ^ iccm_dma_rtag_temp; // @[lib.scala 453:21]
  wire  _T_3161 = |_T_3160; // @[lib.scala 453:29]
  wire [1:0] _T_3165 = io_dma_mem_ctl_dma_mem_addr[3:2] ^ dma_mem_addr_ff; // @[lib.scala 453:21]
  wire  _T_3166 = |_T_3165; // @[lib.scala 453:29]
  wire  _T_3168 = _T_2764 ^ iccm_dma_rvalid_in; // @[lib.scala 475:21]
  wire  _T_3169 = |_T_3168; // @[lib.scala 475:29]
  reg  iccm_dma_rvalid_temp; // @[Reg.scala 27:20]
  wire  _T_3171 = iccm_dma_rvalid_in ^ iccm_dma_rvalid_temp; // @[lib.scala 475:21]
  wire  _T_3172 = |_T_3171; // @[lib.scala 475:29]
  reg  iccm_dma_ecc_error; // @[Reg.scala 27:20]
  wire  _T_3175 = _T_3154 ^ iccm_dma_ecc_error; // @[lib.scala 475:21]
  wire  _T_3176 = |_T_3175; // @[lib.scala 475:29]
  reg [63:0] iccm_dma_rdata_temp; // @[Reg.scala 27:20]
  wire  _T_3180 = _T_2759 & _T_2740; // @[ifu_mem_ctl.scala 558:71]
  wire  _T_3184 = _T_3141 & iccm_correct_ecc; // @[ifu_mem_ctl.scala 559:56]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3185 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [14:0] _T_3187 = _T_3184 ? _T_3185 : io_ifc_fetch_addr_bf[14:0]; // @[ifu_mem_ctl.scala 559:8]
  wire  _T_3579 = _T_3417 == 7'h40; // @[lib.scala 205:62]
  wire  _T_3580 = _T_3567[38] ^ _T_3579; // @[lib.scala 205:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3580,_T_3567[31],_T_3567[15],_T_3567[7],_T_3567[3],_T_3567[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3964 = _T_3802 == 7'h40; // @[lib.scala 205:62]
  wire  _T_3965 = _T_3952[38] ^ _T_3964; // @[lib.scala 205:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3965,_T_3952[31],_T_3952[15],_T_3952[7],_T_3952[3],_T_3952[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3981 = _T_6 & ifc_iccm_access_f; // @[ifu_mem_ctl.scala 571:77]
  wire [1:0] _T_3987 = {iccm_double_ecc_error[0],iccm_double_ecc_error[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_3989 = ifc_iccm_access_f ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_3990 = _T_3987 & _T_3989; // @[ifu_mem_ctl.scala 572:124]
  wire [1:0] _T_3993 = {iccm_double_ecc_error[1],iccm_double_ecc_error[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_3996 = _T_3993 & _T_3989; // @[ifu_mem_ctl.scala 573:66]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[ifu_mem_ctl.scala 580:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[ifu_mem_ctl.scala 581:37]
  reg  iccm_rd_ecc_single_err_ff; // @[Reg.scala 27:20]
  wire  _T_4009 = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[ifu_mem_ctl.scala 585:81]
  wire  iccm_rd_ecc_single_err_hold_in = _T_4009 & _T_339; // @[ifu_mem_ctl.scala 585:110]
  wire  _T_4002 = iccm_rd_ecc_single_err_hold_in ^ iccm_rd_ecc_single_err_ff; // @[lib.scala 475:21]
  wire  _T_4003 = |_T_4002; // @[lib.scala 475:29]
  wire  _T_4005 = ~iccm_rd_ecc_single_err_ff; // @[ifu_mem_ctl.scala 584:93]
  wire  _T_4006 = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err & _T_4005; // @[ifu_mem_ctl.scala 584:91]
  wire  _T_4008 = _T_4006 & _T_339; // @[ifu_mem_ctl.scala 584:121]
  wire  iccm_ecc_write_status = _T_4008 | io_iccm_dma_sb_error; // @[ifu_mem_ctl.scala 584:144]
  reg [13:0] iccm_rw_addr_f; // @[Reg.scala 27:20]
  wire [13:0] _T_4015 = iccm_rw_addr_f + 14'h1; // @[ifu_mem_ctl.scala 588:102]
  wire [13:0] _T_4018 = io_iccm_rw_addr[14:1] ^ iccm_rw_addr_f; // @[lib.scala 453:21]
  wire  _T_4019 = |_T_4018; // @[lib.scala 453:29]
  wire [38:0] _T_4021 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_4026 = ~io_ifc_fetch_uncacheable_bf; // @[ifu_mem_ctl.scala 592:41]
  wire  _T_4027 = io_ifc_fetch_req_bf & _T_4026; // @[ifu_mem_ctl.scala 592:39]
  wire  _T_4029 = _T_4027 & _T_10655; // @[ifu_mem_ctl.scala 592:70]
  wire  _T_4031 = ~miss_state_en; // @[ifu_mem_ctl.scala 593:34]
  wire  _T_4032 = _T_2274 & _T_4031; // @[ifu_mem_ctl.scala 593:32]
  wire  _T_4035 = _T_2290 & _T_4031; // @[ifu_mem_ctl.scala 594:37]
  wire  _T_4036 = _T_4032 | _T_4035; // @[ifu_mem_ctl.scala 593:88]
  wire  _T_4037 = miss_state == 3'h7; // @[ifu_mem_ctl.scala 595:19]
  wire  _T_4039 = _T_4037 & _T_4031; // @[ifu_mem_ctl.scala 595:41]
  wire  _T_4040 = _T_4036 | _T_4039; // @[ifu_mem_ctl.scala 594:88]
  wire  _T_4043 = _T_1281 & _T_4031; // @[ifu_mem_ctl.scala 596:35]
  wire  _T_4044 = _T_4040 | _T_4043; // @[ifu_mem_ctl.scala 595:88]
  wire  _T_4047 = _T_2289 & _T_4031; // @[ifu_mem_ctl.scala 597:38]
  wire  _T_4048 = _T_4044 | _T_4047; // @[ifu_mem_ctl.scala 596:88]
  wire  _T_4050 = _T_2290 & miss_state_en; // @[ifu_mem_ctl.scala 598:37]
  wire  _T_4051 = miss_nxtstate == 3'h3; // @[ifu_mem_ctl.scala 598:71]
  wire  _T_4052 = _T_4050 & _T_4051; // @[ifu_mem_ctl.scala 598:54]
  wire  _T_4053 = _T_4048 | _T_4052; // @[ifu_mem_ctl.scala 597:57]
  wire  _T_4054 = ~_T_4053; // @[ifu_mem_ctl.scala 593:5]
  wire  _T_4055 = _T_4029 & _T_4054; // @[ifu_mem_ctl.scala 592:96]
  wire  _T_4056 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[ifu_mem_ctl.scala 599:26]
  wire  _T_4058 = _T_4056 & _T_4026; // @[ifu_mem_ctl.scala 599:48]
  wire  _T_4060 = _T_4058 & _T_10655; // @[ifu_mem_ctl.scala 599:79]
  wire [1:0] _T_4063 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10530 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[ifu_mem_ctl.scala 687:89]
  wire  bus_wren_1 = _T_10530 & miss_pending; // @[ifu_mem_ctl.scala 687:113]
  wire  _T_10529 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[ifu_mem_ctl.scala 687:89]
  wire  bus_wren_0 = _T_10529 & miss_pending; // @[ifu_mem_ctl.scala 687:113]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_4069 = ~_T_111; // @[ifu_mem_ctl.scala 602:106]
  wire  _T_4070 = _T_2274 & _T_4069; // @[ifu_mem_ctl.scala 602:104]
  wire  _T_4071 = _T_2290 | _T_4070; // @[ifu_mem_ctl.scala 602:77]
  wire  _T_4075 = ~_T_54; // @[ifu_mem_ctl.scala 602:172]
  wire  _T_4076 = _T_4071 & _T_4075; // @[ifu_mem_ctl.scala 602:170]
  wire  _T_4077 = ~_T_4076; // @[ifu_mem_ctl.scala 602:44]
  wire  _T_4080 = io_dec_mem_ctrl_dec_tlu_fence_i_wb ^ reset_all_tags; // @[lib.scala 475:21]
  wire  _T_4081 = |_T_4080; // @[lib.scala 475:29]
  wire  _T_4084 = reset_ic_in | reset_ic_ff; // @[ifu_mem_ctl.scala 605:62]
  wire  _T_4085 = ~_T_4084; // @[ifu_mem_ctl.scala 605:48]
  wire  _T_4086 = _T_282 & _T_4085; // @[ifu_mem_ctl.scala 605:46]
  wire  _T_4087 = ~reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 605:79]
  wire  ic_valid = _T_4086 & _T_4087; // @[ifu_mem_ctl.scala 605:77]
  wire  _T_4089 = debug_c1_clken & io_ic_debug_tag_array; // @[ifu_mem_ctl.scala 606:80]
  wire [6:0] ifu_status_wr_addr_w_debug = _T_4089 ? io_ic_debug_addr[9:3] : ifu_status_wr_addr[11:5]; // @[ifu_mem_ctl.scala 606:39]
  reg [6:0] ifu_status_wr_addr_ff; // @[Reg.scala 27:20]
  wire [6:0] _T_4092 = ifu_status_wr_addr_w_debug ^ ifu_status_wr_addr_ff; // @[lib.scala 453:21]
  wire  _T_4093 = |_T_4092; // @[lib.scala 453:29]
  wire  _T_4095 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[ifu_mem_ctl.scala 611:72]
  wire  _T_10527 = bus_ifu_wr_en_ff_q & last_beat; // @[ifu_mem_ctl.scala 686:43]
  wire  way_status_wr_en = _T_10527 | ic_act_hit_f; // @[ifu_mem_ctl.scala 686:56]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_4095; // @[ifu_mem_ctl.scala 611:51]
  reg  way_status_wr_en_ff; // @[Reg.scala 27:20]
  wire  _T_4096 = way_status_wr_en_w_debug ^ way_status_wr_en_ff; // @[lib.scala 475:21]
  wire  _T_4097 = |_T_4096; // @[lib.scala 475:29]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[ifu_mem_ctl.scala 682:39]
  wire  way_status_new = _T_10527 ? replace_way_mb_any_0 : way_status_hit_new; // @[ifu_mem_ctl.scala 685:24]
  wire  way_status_new_w_debug = _T_4095 ? io_ic_debug_wr_data[4] : way_status_new; // @[ifu_mem_ctl.scala 615:35]
  reg  way_status_new_ff; // @[Reg.scala 27:20]
  wire  _T_4101 = way_status_new_w_debug ^ way_status_new_ff; // @[lib.scala 453:21]
  wire  _T_4102 = |_T_4101; // @[lib.scala 453:29]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[ifu_mem_ctl.scala 619:130]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[ifu_mem_ctl.scala 619:130]
  wire  _T_4121 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[ifu_mem_ctl.scala 623:93]
  wire  _T_4122 = _T_4121 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 623:101]
  wire  _T_4123 = way_status_clken_0 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4126 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[ifu_mem_ctl.scala 623:93]
  wire  _T_4127 = _T_4126 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 623:101]
  wire  _T_4128 = way_status_clken_0 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4131 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[ifu_mem_ctl.scala 623:93]
  wire  _T_4132 = _T_4131 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 623:101]
  wire  _T_4133 = way_status_clken_0 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4136 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[ifu_mem_ctl.scala 623:93]
  wire  _T_4137 = _T_4136 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 623:101]
  wire  _T_4138 = way_status_clken_0 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4141 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[ifu_mem_ctl.scala 623:93]
  wire  _T_4142 = _T_4141 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 623:101]
  wire  _T_4143 = way_status_clken_0 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4146 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[ifu_mem_ctl.scala 623:93]
  wire  _T_4147 = _T_4146 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 623:101]
  wire  _T_4148 = way_status_clken_0 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4151 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[ifu_mem_ctl.scala 623:93]
  wire  _T_4152 = _T_4151 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 623:101]
  wire  _T_4153 = way_status_clken_0 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4156 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[ifu_mem_ctl.scala 623:93]
  wire  _T_4157 = _T_4156 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 623:101]
  wire  _T_4158 = way_status_clken_0 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4163 = way_status_clken_1 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4168 = way_status_clken_1 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4173 = way_status_clken_1 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4178 = way_status_clken_1 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4183 = way_status_clken_1 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4188 = way_status_clken_1 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4193 = way_status_clken_1 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4198 = way_status_clken_1 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4203 = way_status_clken_2 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4208 = way_status_clken_2 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4213 = way_status_clken_2 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4218 = way_status_clken_2 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4223 = way_status_clken_2 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4228 = way_status_clken_2 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4233 = way_status_clken_2 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4238 = way_status_clken_2 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4243 = way_status_clken_3 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4248 = way_status_clken_3 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4253 = way_status_clken_3 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4258 = way_status_clken_3 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4263 = way_status_clken_3 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4268 = way_status_clken_3 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4273 = way_status_clken_3 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4278 = way_status_clken_3 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4283 = way_status_clken_4 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4288 = way_status_clken_4 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4293 = way_status_clken_4 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4298 = way_status_clken_4 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4303 = way_status_clken_4 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4308 = way_status_clken_4 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4313 = way_status_clken_4 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4318 = way_status_clken_4 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4323 = way_status_clken_5 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4328 = way_status_clken_5 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4333 = way_status_clken_5 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4338 = way_status_clken_5 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4343 = way_status_clken_5 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4348 = way_status_clken_5 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4353 = way_status_clken_5 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4358 = way_status_clken_5 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4363 = way_status_clken_6 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4368 = way_status_clken_6 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4373 = way_status_clken_6 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4378 = way_status_clken_6 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4383 = way_status_clken_6 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4388 = way_status_clken_6 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4393 = way_status_clken_6 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4398 = way_status_clken_6 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4403 = way_status_clken_7 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4408 = way_status_clken_7 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4413 = way_status_clken_7 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4418 = way_status_clken_7 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4423 = way_status_clken_7 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4428 = way_status_clken_7 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4433 = way_status_clken_7 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4438 = way_status_clken_7 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4443 = way_status_clken_8 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4448 = way_status_clken_8 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4453 = way_status_clken_8 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4458 = way_status_clken_8 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4463 = way_status_clken_8 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4468 = way_status_clken_8 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4473 = way_status_clken_8 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4478 = way_status_clken_8 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4483 = way_status_clken_9 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4488 = way_status_clken_9 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4493 = way_status_clken_9 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4498 = way_status_clken_9 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4503 = way_status_clken_9 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4508 = way_status_clken_9 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4513 = way_status_clken_9 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4518 = way_status_clken_9 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4523 = way_status_clken_10 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4528 = way_status_clken_10 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4533 = way_status_clken_10 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4538 = way_status_clken_10 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4543 = way_status_clken_10 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4548 = way_status_clken_10 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4553 = way_status_clken_10 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4558 = way_status_clken_10 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4563 = way_status_clken_11 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4568 = way_status_clken_11 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4573 = way_status_clken_11 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4578 = way_status_clken_11 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4583 = way_status_clken_11 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4588 = way_status_clken_11 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4593 = way_status_clken_11 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4598 = way_status_clken_11 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4603 = way_status_clken_12 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4608 = way_status_clken_12 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4613 = way_status_clken_12 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4618 = way_status_clken_12 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4623 = way_status_clken_12 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4628 = way_status_clken_12 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4633 = way_status_clken_12 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4638 = way_status_clken_12 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4643 = way_status_clken_13 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4648 = way_status_clken_13 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4653 = way_status_clken_13 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4658 = way_status_clken_13 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4663 = way_status_clken_13 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4668 = way_status_clken_13 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4673 = way_status_clken_13 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4678 = way_status_clken_13 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4683 = way_status_clken_14 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4688 = way_status_clken_14 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4693 = way_status_clken_14 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4698 = way_status_clken_14 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4703 = way_status_clken_14 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4708 = way_status_clken_14 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4713 = way_status_clken_14 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4718 = way_status_clken_14 & _T_4157; // @[lib.scala 393:57]
  wire  _T_4723 = way_status_clken_15 & _T_4122; // @[lib.scala 393:57]
  wire  _T_4728 = way_status_clken_15 & _T_4127; // @[lib.scala 393:57]
  wire  _T_4733 = way_status_clken_15 & _T_4132; // @[lib.scala 393:57]
  wire  _T_4738 = way_status_clken_15 & _T_4137; // @[lib.scala 393:57]
  wire  _T_4743 = way_status_clken_15 & _T_4142; // @[lib.scala 393:57]
  wire  _T_4748 = way_status_clken_15 & _T_4147; // @[lib.scala 393:57]
  wire  _T_4753 = way_status_clken_15 & _T_4152; // @[lib.scala 393:57]
  wire  _T_4758 = way_status_clken_15 & _T_4157; // @[lib.scala 393:57]
  wire [6:0] ifu_ic_rw_int_addr_w_debug = _T_4089 ? io_ic_debug_addr[9:3] : io_ic_rw_addr[11:5]; // @[ifu_mem_ctl.scala 629:39]
  wire [6:0] _T_5289 = ifu_ic_rw_int_addr_w_debug ^ ifu_ic_rw_int_addr_ff; // @[lib.scala 453:21]
  wire  _T_5290 = |_T_5289; // @[lib.scala 453:29]
  wire  _T_10533 = _T_103 & replace_way_mb_any_1; // @[ifu_mem_ctl.scala 689:82]
  wire  _T_10534 = _T_10533 & miss_pending; // @[ifu_mem_ctl.scala 689:106]
  wire  bus_wren_last_1 = _T_10534 & bus_last_data_beat; // @[ifu_mem_ctl.scala 689:121]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 690:82]
  wire  _T_10536 = bus_wren_last_1 | wren_reset_miss_1; // @[ifu_mem_ctl.scala 691:71]
  wire  _T_10531 = _T_103 & replace_way_mb_any_0; // @[ifu_mem_ctl.scala 689:82]
  wire  _T_10532 = _T_10531 & miss_pending; // @[ifu_mem_ctl.scala 689:106]
  wire  bus_wren_last_0 = _T_10532 & bus_last_data_beat; // @[ifu_mem_ctl.scala 689:121]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 690:82]
  wire  _T_10535 = bus_wren_last_0 | wren_reset_miss_0; // @[ifu_mem_ctl.scala 691:71]
  wire [1:0] ifu_tag_wren = {_T_10536,_T_10535}; // @[Cat.scala 29:58]
  wire [1:0] _T_10587 = _T_4095 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10587 & io_ic_debug_way; // @[ifu_mem_ctl.scala 720:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[ifu_mem_ctl.scala 637:43]
  reg [1:0] ifu_tag_wren_ff; // @[Reg.scala 27:20]
  wire [1:0] _T_5292 = ifu_tag_wren_w_debug ^ ifu_tag_wren_ff; // @[lib.scala 453:21]
  wire  _T_5293 = |_T_5292; // @[lib.scala 453:29]
  wire  ic_valid_w_debug = _T_4095 ? io_ic_debug_wr_data[0] : ic_valid; // @[ifu_mem_ctl.scala 640:29]
  reg  ic_valid_ff; // @[Reg.scala 27:20]
  wire  _T_5297 = ic_valid_w_debug ^ ic_valid_ff; // @[lib.scala 475:21]
  wire  _T_5298 = |_T_5297; // @[lib.scala 475:29]
  wire  _T_5301 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[ifu_mem_ctl.scala 645:76]
  wire  _T_5303 = _T_5301 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 645:85]
  wire  _T_5305 = perr_ic_index_ff[6:5] == 2'h0; // @[ifu_mem_ctl.scala 646:68]
  wire  _T_5307 = _T_5305 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 646:77]
  wire  _T_5308 = _T_5303 | _T_5307; // @[ifu_mem_ctl.scala 645:107]
  wire  _T_5309 = _T_5308 | reset_all_tags; // @[ifu_mem_ctl.scala 646:100]
  wire  _T_5313 = _T_5301 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 645:85]
  wire  _T_5317 = _T_5305 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 646:77]
  wire  _T_5318 = _T_5313 | _T_5317; // @[ifu_mem_ctl.scala 645:107]
  wire  _T_5319 = _T_5318 | reset_all_tags; // @[ifu_mem_ctl.scala 646:100]
  wire [1:0] tag_valid_clken_0 = {_T_5319,_T_5309}; // @[Cat.scala 29:58]
  wire  _T_5321 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[ifu_mem_ctl.scala 645:76]
  wire  _T_5323 = _T_5321 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 645:85]
  wire  _T_5325 = perr_ic_index_ff[6:5] == 2'h1; // @[ifu_mem_ctl.scala 646:68]
  wire  _T_5327 = _T_5325 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 646:77]
  wire  _T_5328 = _T_5323 | _T_5327; // @[ifu_mem_ctl.scala 645:107]
  wire  _T_5329 = _T_5328 | reset_all_tags; // @[ifu_mem_ctl.scala 646:100]
  wire  _T_5333 = _T_5321 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 645:85]
  wire  _T_5337 = _T_5325 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 646:77]
  wire  _T_5338 = _T_5333 | _T_5337; // @[ifu_mem_ctl.scala 645:107]
  wire  _T_5339 = _T_5338 | reset_all_tags; // @[ifu_mem_ctl.scala 646:100]
  wire [1:0] tag_valid_clken_1 = {_T_5339,_T_5329}; // @[Cat.scala 29:58]
  wire  _T_5341 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[ifu_mem_ctl.scala 645:76]
  wire  _T_5343 = _T_5341 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 645:85]
  wire  _T_5345 = perr_ic_index_ff[6:5] == 2'h2; // @[ifu_mem_ctl.scala 646:68]
  wire  _T_5347 = _T_5345 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 646:77]
  wire  _T_5348 = _T_5343 | _T_5347; // @[ifu_mem_ctl.scala 645:107]
  wire  _T_5349 = _T_5348 | reset_all_tags; // @[ifu_mem_ctl.scala 646:100]
  wire  _T_5353 = _T_5341 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 645:85]
  wire  _T_5357 = _T_5345 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 646:77]
  wire  _T_5358 = _T_5353 | _T_5357; // @[ifu_mem_ctl.scala 645:107]
  wire  _T_5359 = _T_5358 | reset_all_tags; // @[ifu_mem_ctl.scala 646:100]
  wire [1:0] tag_valid_clken_2 = {_T_5359,_T_5349}; // @[Cat.scala 29:58]
  wire  _T_5361 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[ifu_mem_ctl.scala 645:76]
  wire  _T_5363 = _T_5361 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 645:85]
  wire  _T_5365 = perr_ic_index_ff[6:5] == 2'h3; // @[ifu_mem_ctl.scala 646:68]
  wire  _T_5367 = _T_5365 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 646:77]
  wire  _T_5368 = _T_5363 | _T_5367; // @[ifu_mem_ctl.scala 645:107]
  wire  _T_5369 = _T_5368 | reset_all_tags; // @[ifu_mem_ctl.scala 646:100]
  wire  _T_5373 = _T_5361 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 645:85]
  wire  _T_5377 = _T_5365 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 646:77]
  wire  _T_5378 = _T_5373 | _T_5377; // @[ifu_mem_ctl.scala 645:107]
  wire  _T_5379 = _T_5378 | reset_all_tags; // @[ifu_mem_ctl.scala 646:100]
  wire [1:0] tag_valid_clken_3 = {_T_5379,_T_5369}; // @[Cat.scala 29:58]
  wire  _T_5390 = ic_valid_ff & _T_198; // @[ifu_mem_ctl.scala 654:66]
  wire  _T_5391 = ~perr_sel_invalidate; // @[ifu_mem_ctl.scala 654:93]
  wire  _T_5392 = _T_5390 & _T_5391; // @[ifu_mem_ctl.scala 654:91]
  wire  _T_5395 = _T_4900 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5396 = perr_ic_index_ff == 7'h0; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5398 = _T_5396 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5399 = _T_5395 | _T_5398; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5400 = _T_5399 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5403 = tag_valid_clken_0[0] & _T_5400; // @[lib.scala 393:57]
  wire  _T_5412 = _T_4901 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5413 = perr_ic_index_ff == 7'h1; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5415 = _T_5413 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5416 = _T_5412 | _T_5415; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5417 = _T_5416 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5420 = tag_valid_clken_0[0] & _T_5417; // @[lib.scala 393:57]
  wire  _T_5429 = _T_4902 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5430 = perr_ic_index_ff == 7'h2; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5432 = _T_5430 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5433 = _T_5429 | _T_5432; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5434 = _T_5433 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5437 = tag_valid_clken_0[0] & _T_5434; // @[lib.scala 393:57]
  wire  _T_5446 = _T_4903 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5447 = perr_ic_index_ff == 7'h3; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5449 = _T_5447 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5450 = _T_5446 | _T_5449; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5451 = _T_5450 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5454 = tag_valid_clken_0[0] & _T_5451; // @[lib.scala 393:57]
  wire  _T_5463 = _T_4904 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5464 = perr_ic_index_ff == 7'h4; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5466 = _T_5464 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5467 = _T_5463 | _T_5466; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5468 = _T_5467 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5471 = tag_valid_clken_0[0] & _T_5468; // @[lib.scala 393:57]
  wire  _T_5480 = _T_4905 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5481 = perr_ic_index_ff == 7'h5; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5483 = _T_5481 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5484 = _T_5480 | _T_5483; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5485 = _T_5484 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5488 = tag_valid_clken_0[0] & _T_5485; // @[lib.scala 393:57]
  wire  _T_5497 = _T_4906 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5498 = perr_ic_index_ff == 7'h6; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5500 = _T_5498 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5501 = _T_5497 | _T_5500; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5502 = _T_5501 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5505 = tag_valid_clken_0[0] & _T_5502; // @[lib.scala 393:57]
  wire  _T_5514 = _T_4907 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5515 = perr_ic_index_ff == 7'h7; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5517 = _T_5515 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5518 = _T_5514 | _T_5517; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5519 = _T_5518 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5522 = tag_valid_clken_0[0] & _T_5519; // @[lib.scala 393:57]
  wire  _T_5531 = _T_4908 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5532 = perr_ic_index_ff == 7'h8; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5534 = _T_5532 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5535 = _T_5531 | _T_5534; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5536 = _T_5535 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5539 = tag_valid_clken_0[0] & _T_5536; // @[lib.scala 393:57]
  wire  _T_5548 = _T_4909 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5549 = perr_ic_index_ff == 7'h9; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5551 = _T_5549 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5552 = _T_5548 | _T_5551; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5553 = _T_5552 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5556 = tag_valid_clken_0[0] & _T_5553; // @[lib.scala 393:57]
  wire  _T_5565 = _T_4910 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5566 = perr_ic_index_ff == 7'ha; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5568 = _T_5566 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5569 = _T_5565 | _T_5568; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5570 = _T_5569 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5573 = tag_valid_clken_0[0] & _T_5570; // @[lib.scala 393:57]
  wire  _T_5582 = _T_4911 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5583 = perr_ic_index_ff == 7'hb; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5585 = _T_5583 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5586 = _T_5582 | _T_5585; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5587 = _T_5586 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5590 = tag_valid_clken_0[0] & _T_5587; // @[lib.scala 393:57]
  wire  _T_5599 = _T_4912 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5600 = perr_ic_index_ff == 7'hc; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5602 = _T_5600 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5603 = _T_5599 | _T_5602; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5604 = _T_5603 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5607 = tag_valid_clken_0[0] & _T_5604; // @[lib.scala 393:57]
  wire  _T_5616 = _T_4913 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5617 = perr_ic_index_ff == 7'hd; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5619 = _T_5617 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5620 = _T_5616 | _T_5619; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5621 = _T_5620 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5624 = tag_valid_clken_0[0] & _T_5621; // @[lib.scala 393:57]
  wire  _T_5633 = _T_4914 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5634 = perr_ic_index_ff == 7'he; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5636 = _T_5634 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5637 = _T_5633 | _T_5636; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5638 = _T_5637 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5641 = tag_valid_clken_0[0] & _T_5638; // @[lib.scala 393:57]
  wire  _T_5650 = _T_4915 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5651 = perr_ic_index_ff == 7'hf; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5653 = _T_5651 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5654 = _T_5650 | _T_5653; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5655 = _T_5654 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5658 = tag_valid_clken_0[0] & _T_5655; // @[lib.scala 393:57]
  wire  _T_5667 = _T_4916 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5668 = perr_ic_index_ff == 7'h10; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5670 = _T_5668 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5671 = _T_5667 | _T_5670; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5672 = _T_5671 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5675 = tag_valid_clken_0[0] & _T_5672; // @[lib.scala 393:57]
  wire  _T_5684 = _T_4917 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5685 = perr_ic_index_ff == 7'h11; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5687 = _T_5685 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5688 = _T_5684 | _T_5687; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5689 = _T_5688 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5692 = tag_valid_clken_0[0] & _T_5689; // @[lib.scala 393:57]
  wire  _T_5701 = _T_4918 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5702 = perr_ic_index_ff == 7'h12; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5704 = _T_5702 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5705 = _T_5701 | _T_5704; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5706 = _T_5705 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5709 = tag_valid_clken_0[0] & _T_5706; // @[lib.scala 393:57]
  wire  _T_5718 = _T_4919 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5719 = perr_ic_index_ff == 7'h13; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5721 = _T_5719 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5722 = _T_5718 | _T_5721; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5723 = _T_5722 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5726 = tag_valid_clken_0[0] & _T_5723; // @[lib.scala 393:57]
  wire  _T_5735 = _T_4920 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5736 = perr_ic_index_ff == 7'h14; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5738 = _T_5736 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5739 = _T_5735 | _T_5738; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5740 = _T_5739 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5743 = tag_valid_clken_0[0] & _T_5740; // @[lib.scala 393:57]
  wire  _T_5752 = _T_4921 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5753 = perr_ic_index_ff == 7'h15; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5755 = _T_5753 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5756 = _T_5752 | _T_5755; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5757 = _T_5756 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5760 = tag_valid_clken_0[0] & _T_5757; // @[lib.scala 393:57]
  wire  _T_5769 = _T_4922 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5770 = perr_ic_index_ff == 7'h16; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5772 = _T_5770 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5773 = _T_5769 | _T_5772; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5774 = _T_5773 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5777 = tag_valid_clken_0[0] & _T_5774; // @[lib.scala 393:57]
  wire  _T_5786 = _T_4923 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5787 = perr_ic_index_ff == 7'h17; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5789 = _T_5787 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5790 = _T_5786 | _T_5789; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5791 = _T_5790 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5794 = tag_valid_clken_0[0] & _T_5791; // @[lib.scala 393:57]
  wire  _T_5803 = _T_4924 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5804 = perr_ic_index_ff == 7'h18; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5806 = _T_5804 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5807 = _T_5803 | _T_5806; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5808 = _T_5807 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5811 = tag_valid_clken_0[0] & _T_5808; // @[lib.scala 393:57]
  wire  _T_5820 = _T_4925 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5821 = perr_ic_index_ff == 7'h19; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5823 = _T_5821 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5824 = _T_5820 | _T_5823; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5825 = _T_5824 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5828 = tag_valid_clken_0[0] & _T_5825; // @[lib.scala 393:57]
  wire  _T_5837 = _T_4926 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5838 = perr_ic_index_ff == 7'h1a; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5840 = _T_5838 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5841 = _T_5837 | _T_5840; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5842 = _T_5841 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5845 = tag_valid_clken_0[0] & _T_5842; // @[lib.scala 393:57]
  wire  _T_5854 = _T_4927 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5855 = perr_ic_index_ff == 7'h1b; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5857 = _T_5855 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5858 = _T_5854 | _T_5857; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5859 = _T_5858 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5862 = tag_valid_clken_0[0] & _T_5859; // @[lib.scala 393:57]
  wire  _T_5871 = _T_4928 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5872 = perr_ic_index_ff == 7'h1c; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5874 = _T_5872 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5875 = _T_5871 | _T_5874; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5876 = _T_5875 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5879 = tag_valid_clken_0[0] & _T_5876; // @[lib.scala 393:57]
  wire  _T_5888 = _T_4929 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5889 = perr_ic_index_ff == 7'h1d; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5891 = _T_5889 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5892 = _T_5888 | _T_5891; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5893 = _T_5892 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5896 = tag_valid_clken_0[0] & _T_5893; // @[lib.scala 393:57]
  wire  _T_5905 = _T_4930 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5906 = perr_ic_index_ff == 7'h1e; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5908 = _T_5906 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5909 = _T_5905 | _T_5908; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5910 = _T_5909 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5913 = tag_valid_clken_0[0] & _T_5910; // @[lib.scala 393:57]
  wire  _T_5922 = _T_4931 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5923 = perr_ic_index_ff == 7'h1f; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_5925 = _T_5923 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5926 = _T_5922 | _T_5925; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5927 = _T_5926 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5930 = tag_valid_clken_0[0] & _T_5927; // @[lib.scala 393:57]
  wire  _T_5939 = _T_4900 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5942 = _T_5396 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5943 = _T_5939 | _T_5942; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5944 = _T_5943 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5947 = tag_valid_clken_0[1] & _T_5944; // @[lib.scala 393:57]
  wire  _T_5956 = _T_4901 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5959 = _T_5413 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5960 = _T_5956 | _T_5959; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5961 = _T_5960 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5964 = tag_valid_clken_0[1] & _T_5961; // @[lib.scala 393:57]
  wire  _T_5973 = _T_4902 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5976 = _T_5430 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5977 = _T_5973 | _T_5976; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5978 = _T_5977 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5981 = tag_valid_clken_0[1] & _T_5978; // @[lib.scala 393:57]
  wire  _T_5990 = _T_4903 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_5993 = _T_5447 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_5994 = _T_5990 | _T_5993; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_5995 = _T_5994 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_5998 = tag_valid_clken_0[1] & _T_5995; // @[lib.scala 393:57]
  wire  _T_6007 = _T_4904 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6010 = _T_5464 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6011 = _T_6007 | _T_6010; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6012 = _T_6011 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6015 = tag_valid_clken_0[1] & _T_6012; // @[lib.scala 393:57]
  wire  _T_6024 = _T_4905 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6027 = _T_5481 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6028 = _T_6024 | _T_6027; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6029 = _T_6028 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6032 = tag_valid_clken_0[1] & _T_6029; // @[lib.scala 393:57]
  wire  _T_6041 = _T_4906 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6044 = _T_5498 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6045 = _T_6041 | _T_6044; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6046 = _T_6045 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6049 = tag_valid_clken_0[1] & _T_6046; // @[lib.scala 393:57]
  wire  _T_6058 = _T_4907 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6061 = _T_5515 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6062 = _T_6058 | _T_6061; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6063 = _T_6062 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6066 = tag_valid_clken_0[1] & _T_6063; // @[lib.scala 393:57]
  wire  _T_6075 = _T_4908 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6078 = _T_5532 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6079 = _T_6075 | _T_6078; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6080 = _T_6079 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6083 = tag_valid_clken_0[1] & _T_6080; // @[lib.scala 393:57]
  wire  _T_6092 = _T_4909 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6095 = _T_5549 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6096 = _T_6092 | _T_6095; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6097 = _T_6096 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6100 = tag_valid_clken_0[1] & _T_6097; // @[lib.scala 393:57]
  wire  _T_6109 = _T_4910 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6112 = _T_5566 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6113 = _T_6109 | _T_6112; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6114 = _T_6113 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6117 = tag_valid_clken_0[1] & _T_6114; // @[lib.scala 393:57]
  wire  _T_6126 = _T_4911 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6129 = _T_5583 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6130 = _T_6126 | _T_6129; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6131 = _T_6130 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6134 = tag_valid_clken_0[1] & _T_6131; // @[lib.scala 393:57]
  wire  _T_6143 = _T_4912 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6146 = _T_5600 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6147 = _T_6143 | _T_6146; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6148 = _T_6147 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6151 = tag_valid_clken_0[1] & _T_6148; // @[lib.scala 393:57]
  wire  _T_6160 = _T_4913 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6163 = _T_5617 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6164 = _T_6160 | _T_6163; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6165 = _T_6164 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6168 = tag_valid_clken_0[1] & _T_6165; // @[lib.scala 393:57]
  wire  _T_6177 = _T_4914 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6180 = _T_5634 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6181 = _T_6177 | _T_6180; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6182 = _T_6181 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6185 = tag_valid_clken_0[1] & _T_6182; // @[lib.scala 393:57]
  wire  _T_6194 = _T_4915 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6197 = _T_5651 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6198 = _T_6194 | _T_6197; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6199 = _T_6198 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6202 = tag_valid_clken_0[1] & _T_6199; // @[lib.scala 393:57]
  wire  _T_6211 = _T_4916 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6214 = _T_5668 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6215 = _T_6211 | _T_6214; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6216 = _T_6215 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6219 = tag_valid_clken_0[1] & _T_6216; // @[lib.scala 393:57]
  wire  _T_6228 = _T_4917 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6231 = _T_5685 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6232 = _T_6228 | _T_6231; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6233 = _T_6232 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6236 = tag_valid_clken_0[1] & _T_6233; // @[lib.scala 393:57]
  wire  _T_6245 = _T_4918 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6248 = _T_5702 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6249 = _T_6245 | _T_6248; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6250 = _T_6249 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6253 = tag_valid_clken_0[1] & _T_6250; // @[lib.scala 393:57]
  wire  _T_6262 = _T_4919 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6265 = _T_5719 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6266 = _T_6262 | _T_6265; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6267 = _T_6266 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6270 = tag_valid_clken_0[1] & _T_6267; // @[lib.scala 393:57]
  wire  _T_6279 = _T_4920 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6282 = _T_5736 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6283 = _T_6279 | _T_6282; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6284 = _T_6283 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6287 = tag_valid_clken_0[1] & _T_6284; // @[lib.scala 393:57]
  wire  _T_6296 = _T_4921 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6299 = _T_5753 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6300 = _T_6296 | _T_6299; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6301 = _T_6300 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6304 = tag_valid_clken_0[1] & _T_6301; // @[lib.scala 393:57]
  wire  _T_6313 = _T_4922 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6316 = _T_5770 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6317 = _T_6313 | _T_6316; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6318 = _T_6317 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6321 = tag_valid_clken_0[1] & _T_6318; // @[lib.scala 393:57]
  wire  _T_6330 = _T_4923 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6333 = _T_5787 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6334 = _T_6330 | _T_6333; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6335 = _T_6334 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6338 = tag_valid_clken_0[1] & _T_6335; // @[lib.scala 393:57]
  wire  _T_6347 = _T_4924 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6350 = _T_5804 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6351 = _T_6347 | _T_6350; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6352 = _T_6351 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6355 = tag_valid_clken_0[1] & _T_6352; // @[lib.scala 393:57]
  wire  _T_6364 = _T_4925 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6367 = _T_5821 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6368 = _T_6364 | _T_6367; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6369 = _T_6368 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6372 = tag_valid_clken_0[1] & _T_6369; // @[lib.scala 393:57]
  wire  _T_6381 = _T_4926 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6384 = _T_5838 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6385 = _T_6381 | _T_6384; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6386 = _T_6385 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6389 = tag_valid_clken_0[1] & _T_6386; // @[lib.scala 393:57]
  wire  _T_6398 = _T_4927 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6401 = _T_5855 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6402 = _T_6398 | _T_6401; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6403 = _T_6402 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6406 = tag_valid_clken_0[1] & _T_6403; // @[lib.scala 393:57]
  wire  _T_6415 = _T_4928 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6418 = _T_5872 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6419 = _T_6415 | _T_6418; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6420 = _T_6419 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6423 = tag_valid_clken_0[1] & _T_6420; // @[lib.scala 393:57]
  wire  _T_6432 = _T_4929 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6435 = _T_5889 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6436 = _T_6432 | _T_6435; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6437 = _T_6436 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6440 = tag_valid_clken_0[1] & _T_6437; // @[lib.scala 393:57]
  wire  _T_6449 = _T_4930 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6452 = _T_5906 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6453 = _T_6449 | _T_6452; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6454 = _T_6453 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6457 = tag_valid_clken_0[1] & _T_6454; // @[lib.scala 393:57]
  wire  _T_6466 = _T_4931 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6469 = _T_5923 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6470 = _T_6466 | _T_6469; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6471 = _T_6470 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6474 = tag_valid_clken_0[1] & _T_6471; // @[lib.scala 393:57]
  wire  _T_6483 = _T_4932 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6484 = perr_ic_index_ff == 7'h20; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6486 = _T_6484 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6487 = _T_6483 | _T_6486; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6488 = _T_6487 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6491 = tag_valid_clken_1[0] & _T_6488; // @[lib.scala 393:57]
  wire  _T_6500 = _T_4933 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6501 = perr_ic_index_ff == 7'h21; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6503 = _T_6501 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6504 = _T_6500 | _T_6503; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6505 = _T_6504 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6508 = tag_valid_clken_1[0] & _T_6505; // @[lib.scala 393:57]
  wire  _T_6517 = _T_4934 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6518 = perr_ic_index_ff == 7'h22; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6520 = _T_6518 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6521 = _T_6517 | _T_6520; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6522 = _T_6521 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6525 = tag_valid_clken_1[0] & _T_6522; // @[lib.scala 393:57]
  wire  _T_6534 = _T_4935 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6535 = perr_ic_index_ff == 7'h23; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6537 = _T_6535 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6538 = _T_6534 | _T_6537; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6539 = _T_6538 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6542 = tag_valid_clken_1[0] & _T_6539; // @[lib.scala 393:57]
  wire  _T_6551 = _T_4936 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6552 = perr_ic_index_ff == 7'h24; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6554 = _T_6552 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6555 = _T_6551 | _T_6554; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6556 = _T_6555 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6559 = tag_valid_clken_1[0] & _T_6556; // @[lib.scala 393:57]
  wire  _T_6568 = _T_4937 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6569 = perr_ic_index_ff == 7'h25; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6571 = _T_6569 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6572 = _T_6568 | _T_6571; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6573 = _T_6572 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6576 = tag_valid_clken_1[0] & _T_6573; // @[lib.scala 393:57]
  wire  _T_6585 = _T_4938 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6586 = perr_ic_index_ff == 7'h26; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6588 = _T_6586 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6589 = _T_6585 | _T_6588; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6590 = _T_6589 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6593 = tag_valid_clken_1[0] & _T_6590; // @[lib.scala 393:57]
  wire  _T_6602 = _T_4939 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6603 = perr_ic_index_ff == 7'h27; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6605 = _T_6603 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6606 = _T_6602 | _T_6605; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6607 = _T_6606 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6610 = tag_valid_clken_1[0] & _T_6607; // @[lib.scala 393:57]
  wire  _T_6619 = _T_4940 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6620 = perr_ic_index_ff == 7'h28; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6622 = _T_6620 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6623 = _T_6619 | _T_6622; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6624 = _T_6623 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6627 = tag_valid_clken_1[0] & _T_6624; // @[lib.scala 393:57]
  wire  _T_6636 = _T_4941 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6637 = perr_ic_index_ff == 7'h29; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6639 = _T_6637 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6640 = _T_6636 | _T_6639; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6641 = _T_6640 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6644 = tag_valid_clken_1[0] & _T_6641; // @[lib.scala 393:57]
  wire  _T_6653 = _T_4942 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6654 = perr_ic_index_ff == 7'h2a; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6656 = _T_6654 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6657 = _T_6653 | _T_6656; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6658 = _T_6657 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6661 = tag_valid_clken_1[0] & _T_6658; // @[lib.scala 393:57]
  wire  _T_6670 = _T_4943 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6671 = perr_ic_index_ff == 7'h2b; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6673 = _T_6671 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6674 = _T_6670 | _T_6673; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6675 = _T_6674 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6678 = tag_valid_clken_1[0] & _T_6675; // @[lib.scala 393:57]
  wire  _T_6687 = _T_4944 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6688 = perr_ic_index_ff == 7'h2c; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6690 = _T_6688 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6691 = _T_6687 | _T_6690; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6692 = _T_6691 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6695 = tag_valid_clken_1[0] & _T_6692; // @[lib.scala 393:57]
  wire  _T_6704 = _T_4945 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6705 = perr_ic_index_ff == 7'h2d; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6707 = _T_6705 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6708 = _T_6704 | _T_6707; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6709 = _T_6708 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6712 = tag_valid_clken_1[0] & _T_6709; // @[lib.scala 393:57]
  wire  _T_6721 = _T_4946 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6722 = perr_ic_index_ff == 7'h2e; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6724 = _T_6722 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6725 = _T_6721 | _T_6724; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6726 = _T_6725 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6729 = tag_valid_clken_1[0] & _T_6726; // @[lib.scala 393:57]
  wire  _T_6738 = _T_4947 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6739 = perr_ic_index_ff == 7'h2f; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6741 = _T_6739 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6742 = _T_6738 | _T_6741; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6743 = _T_6742 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6746 = tag_valid_clken_1[0] & _T_6743; // @[lib.scala 393:57]
  wire  _T_6755 = _T_4948 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6756 = perr_ic_index_ff == 7'h30; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6758 = _T_6756 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6759 = _T_6755 | _T_6758; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6760 = _T_6759 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6763 = tag_valid_clken_1[0] & _T_6760; // @[lib.scala 393:57]
  wire  _T_6772 = _T_4949 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6773 = perr_ic_index_ff == 7'h31; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6775 = _T_6773 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6776 = _T_6772 | _T_6775; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6777 = _T_6776 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6780 = tag_valid_clken_1[0] & _T_6777; // @[lib.scala 393:57]
  wire  _T_6789 = _T_4950 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6790 = perr_ic_index_ff == 7'h32; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6792 = _T_6790 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6793 = _T_6789 | _T_6792; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6794 = _T_6793 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6797 = tag_valid_clken_1[0] & _T_6794; // @[lib.scala 393:57]
  wire  _T_6806 = _T_4951 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6807 = perr_ic_index_ff == 7'h33; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6809 = _T_6807 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6810 = _T_6806 | _T_6809; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6811 = _T_6810 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6814 = tag_valid_clken_1[0] & _T_6811; // @[lib.scala 393:57]
  wire  _T_6823 = _T_4952 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6824 = perr_ic_index_ff == 7'h34; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6826 = _T_6824 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6827 = _T_6823 | _T_6826; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6828 = _T_6827 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6831 = tag_valid_clken_1[0] & _T_6828; // @[lib.scala 393:57]
  wire  _T_6840 = _T_4953 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6841 = perr_ic_index_ff == 7'h35; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6843 = _T_6841 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6844 = _T_6840 | _T_6843; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6845 = _T_6844 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6848 = tag_valid_clken_1[0] & _T_6845; // @[lib.scala 393:57]
  wire  _T_6857 = _T_4954 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6858 = perr_ic_index_ff == 7'h36; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6860 = _T_6858 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6861 = _T_6857 | _T_6860; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6862 = _T_6861 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6865 = tag_valid_clken_1[0] & _T_6862; // @[lib.scala 393:57]
  wire  _T_6874 = _T_4955 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6875 = perr_ic_index_ff == 7'h37; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6877 = _T_6875 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6878 = _T_6874 | _T_6877; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6879 = _T_6878 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6882 = tag_valid_clken_1[0] & _T_6879; // @[lib.scala 393:57]
  wire  _T_6891 = _T_4956 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6892 = perr_ic_index_ff == 7'h38; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6894 = _T_6892 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6895 = _T_6891 | _T_6894; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6896 = _T_6895 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6899 = tag_valid_clken_1[0] & _T_6896; // @[lib.scala 393:57]
  wire  _T_6908 = _T_4957 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6909 = perr_ic_index_ff == 7'h39; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6911 = _T_6909 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6912 = _T_6908 | _T_6911; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6913 = _T_6912 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6916 = tag_valid_clken_1[0] & _T_6913; // @[lib.scala 393:57]
  wire  _T_6925 = _T_4958 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6926 = perr_ic_index_ff == 7'h3a; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6928 = _T_6926 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6929 = _T_6925 | _T_6928; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6930 = _T_6929 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6933 = tag_valid_clken_1[0] & _T_6930; // @[lib.scala 393:57]
  wire  _T_6942 = _T_4959 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6943 = perr_ic_index_ff == 7'h3b; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6945 = _T_6943 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6946 = _T_6942 | _T_6945; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6947 = _T_6946 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6950 = tag_valid_clken_1[0] & _T_6947; // @[lib.scala 393:57]
  wire  _T_6959 = _T_4960 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6960 = perr_ic_index_ff == 7'h3c; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6962 = _T_6960 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6963 = _T_6959 | _T_6962; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6964 = _T_6963 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6967 = tag_valid_clken_1[0] & _T_6964; // @[lib.scala 393:57]
  wire  _T_6976 = _T_4961 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6977 = perr_ic_index_ff == 7'h3d; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6979 = _T_6977 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6980 = _T_6976 | _T_6979; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6981 = _T_6980 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_6984 = tag_valid_clken_1[0] & _T_6981; // @[lib.scala 393:57]
  wire  _T_6993 = _T_4962 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_6994 = perr_ic_index_ff == 7'h3e; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_6996 = _T_6994 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_6997 = _T_6993 | _T_6996; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_6998 = _T_6997 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7001 = tag_valid_clken_1[0] & _T_6998; // @[lib.scala 393:57]
  wire  _T_7010 = _T_4963 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7011 = perr_ic_index_ff == 7'h3f; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7013 = _T_7011 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7014 = _T_7010 | _T_7013; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7015 = _T_7014 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7018 = tag_valid_clken_1[0] & _T_7015; // @[lib.scala 393:57]
  wire  _T_7027 = _T_4932 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7030 = _T_6484 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7031 = _T_7027 | _T_7030; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7032 = _T_7031 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7035 = tag_valid_clken_1[1] & _T_7032; // @[lib.scala 393:57]
  wire  _T_7044 = _T_4933 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7047 = _T_6501 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7048 = _T_7044 | _T_7047; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7049 = _T_7048 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7052 = tag_valid_clken_1[1] & _T_7049; // @[lib.scala 393:57]
  wire  _T_7061 = _T_4934 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7064 = _T_6518 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7065 = _T_7061 | _T_7064; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7066 = _T_7065 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7069 = tag_valid_clken_1[1] & _T_7066; // @[lib.scala 393:57]
  wire  _T_7078 = _T_4935 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7081 = _T_6535 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7082 = _T_7078 | _T_7081; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7083 = _T_7082 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7086 = tag_valid_clken_1[1] & _T_7083; // @[lib.scala 393:57]
  wire  _T_7095 = _T_4936 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7098 = _T_6552 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7099 = _T_7095 | _T_7098; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7100 = _T_7099 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7103 = tag_valid_clken_1[1] & _T_7100; // @[lib.scala 393:57]
  wire  _T_7112 = _T_4937 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7115 = _T_6569 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7116 = _T_7112 | _T_7115; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7117 = _T_7116 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7120 = tag_valid_clken_1[1] & _T_7117; // @[lib.scala 393:57]
  wire  _T_7129 = _T_4938 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7132 = _T_6586 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7133 = _T_7129 | _T_7132; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7134 = _T_7133 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7137 = tag_valid_clken_1[1] & _T_7134; // @[lib.scala 393:57]
  wire  _T_7146 = _T_4939 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7149 = _T_6603 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7150 = _T_7146 | _T_7149; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7151 = _T_7150 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7154 = tag_valid_clken_1[1] & _T_7151; // @[lib.scala 393:57]
  wire  _T_7163 = _T_4940 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7166 = _T_6620 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7167 = _T_7163 | _T_7166; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7168 = _T_7167 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7171 = tag_valid_clken_1[1] & _T_7168; // @[lib.scala 393:57]
  wire  _T_7180 = _T_4941 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7183 = _T_6637 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7184 = _T_7180 | _T_7183; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7185 = _T_7184 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7188 = tag_valid_clken_1[1] & _T_7185; // @[lib.scala 393:57]
  wire  _T_7197 = _T_4942 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7200 = _T_6654 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7201 = _T_7197 | _T_7200; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7202 = _T_7201 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7205 = tag_valid_clken_1[1] & _T_7202; // @[lib.scala 393:57]
  wire  _T_7214 = _T_4943 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7217 = _T_6671 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7218 = _T_7214 | _T_7217; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7219 = _T_7218 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7222 = tag_valid_clken_1[1] & _T_7219; // @[lib.scala 393:57]
  wire  _T_7231 = _T_4944 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7234 = _T_6688 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7235 = _T_7231 | _T_7234; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7236 = _T_7235 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7239 = tag_valid_clken_1[1] & _T_7236; // @[lib.scala 393:57]
  wire  _T_7248 = _T_4945 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7251 = _T_6705 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7252 = _T_7248 | _T_7251; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7253 = _T_7252 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7256 = tag_valid_clken_1[1] & _T_7253; // @[lib.scala 393:57]
  wire  _T_7265 = _T_4946 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7268 = _T_6722 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7269 = _T_7265 | _T_7268; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7270 = _T_7269 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7273 = tag_valid_clken_1[1] & _T_7270; // @[lib.scala 393:57]
  wire  _T_7282 = _T_4947 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7285 = _T_6739 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7286 = _T_7282 | _T_7285; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7287 = _T_7286 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7290 = tag_valid_clken_1[1] & _T_7287; // @[lib.scala 393:57]
  wire  _T_7299 = _T_4948 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7302 = _T_6756 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7303 = _T_7299 | _T_7302; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7304 = _T_7303 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7307 = tag_valid_clken_1[1] & _T_7304; // @[lib.scala 393:57]
  wire  _T_7316 = _T_4949 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7319 = _T_6773 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7320 = _T_7316 | _T_7319; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7321 = _T_7320 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7324 = tag_valid_clken_1[1] & _T_7321; // @[lib.scala 393:57]
  wire  _T_7333 = _T_4950 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7336 = _T_6790 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7337 = _T_7333 | _T_7336; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7338 = _T_7337 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7341 = tag_valid_clken_1[1] & _T_7338; // @[lib.scala 393:57]
  wire  _T_7350 = _T_4951 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7353 = _T_6807 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7354 = _T_7350 | _T_7353; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7355 = _T_7354 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7358 = tag_valid_clken_1[1] & _T_7355; // @[lib.scala 393:57]
  wire  _T_7367 = _T_4952 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7370 = _T_6824 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7371 = _T_7367 | _T_7370; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7372 = _T_7371 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7375 = tag_valid_clken_1[1] & _T_7372; // @[lib.scala 393:57]
  wire  _T_7384 = _T_4953 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7387 = _T_6841 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7388 = _T_7384 | _T_7387; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7389 = _T_7388 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7392 = tag_valid_clken_1[1] & _T_7389; // @[lib.scala 393:57]
  wire  _T_7401 = _T_4954 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7404 = _T_6858 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7405 = _T_7401 | _T_7404; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7406 = _T_7405 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7409 = tag_valid_clken_1[1] & _T_7406; // @[lib.scala 393:57]
  wire  _T_7418 = _T_4955 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7421 = _T_6875 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7422 = _T_7418 | _T_7421; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7423 = _T_7422 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7426 = tag_valid_clken_1[1] & _T_7423; // @[lib.scala 393:57]
  wire  _T_7435 = _T_4956 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7438 = _T_6892 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7439 = _T_7435 | _T_7438; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7440 = _T_7439 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7443 = tag_valid_clken_1[1] & _T_7440; // @[lib.scala 393:57]
  wire  _T_7452 = _T_4957 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7455 = _T_6909 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7456 = _T_7452 | _T_7455; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7457 = _T_7456 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7460 = tag_valid_clken_1[1] & _T_7457; // @[lib.scala 393:57]
  wire  _T_7469 = _T_4958 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7472 = _T_6926 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7473 = _T_7469 | _T_7472; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7474 = _T_7473 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7477 = tag_valid_clken_1[1] & _T_7474; // @[lib.scala 393:57]
  wire  _T_7486 = _T_4959 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7489 = _T_6943 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7490 = _T_7486 | _T_7489; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7491 = _T_7490 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7494 = tag_valid_clken_1[1] & _T_7491; // @[lib.scala 393:57]
  wire  _T_7503 = _T_4960 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7506 = _T_6960 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7507 = _T_7503 | _T_7506; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7508 = _T_7507 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7511 = tag_valid_clken_1[1] & _T_7508; // @[lib.scala 393:57]
  wire  _T_7520 = _T_4961 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7523 = _T_6977 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7524 = _T_7520 | _T_7523; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7525 = _T_7524 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7528 = tag_valid_clken_1[1] & _T_7525; // @[lib.scala 393:57]
  wire  _T_7537 = _T_4962 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7540 = _T_6994 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7541 = _T_7537 | _T_7540; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7542 = _T_7541 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7545 = tag_valid_clken_1[1] & _T_7542; // @[lib.scala 393:57]
  wire  _T_7554 = _T_4963 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7557 = _T_7011 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7558 = _T_7554 | _T_7557; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7559 = _T_7558 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7562 = tag_valid_clken_1[1] & _T_7559; // @[lib.scala 393:57]
  wire  _T_7571 = _T_4964 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7572 = perr_ic_index_ff == 7'h40; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7574 = _T_7572 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7575 = _T_7571 | _T_7574; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7576 = _T_7575 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7579 = tag_valid_clken_2[0] & _T_7576; // @[lib.scala 393:57]
  wire  _T_7588 = _T_4965 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7589 = perr_ic_index_ff == 7'h41; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7591 = _T_7589 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7592 = _T_7588 | _T_7591; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7593 = _T_7592 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7596 = tag_valid_clken_2[0] & _T_7593; // @[lib.scala 393:57]
  wire  _T_7605 = _T_4966 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7606 = perr_ic_index_ff == 7'h42; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7608 = _T_7606 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7609 = _T_7605 | _T_7608; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7610 = _T_7609 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7613 = tag_valid_clken_2[0] & _T_7610; // @[lib.scala 393:57]
  wire  _T_7622 = _T_4967 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7623 = perr_ic_index_ff == 7'h43; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7625 = _T_7623 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7626 = _T_7622 | _T_7625; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7627 = _T_7626 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7630 = tag_valid_clken_2[0] & _T_7627; // @[lib.scala 393:57]
  wire  _T_7639 = _T_4968 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7640 = perr_ic_index_ff == 7'h44; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7642 = _T_7640 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7643 = _T_7639 | _T_7642; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7644 = _T_7643 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7647 = tag_valid_clken_2[0] & _T_7644; // @[lib.scala 393:57]
  wire  _T_7656 = _T_4969 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7657 = perr_ic_index_ff == 7'h45; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7659 = _T_7657 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7660 = _T_7656 | _T_7659; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7661 = _T_7660 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7664 = tag_valid_clken_2[0] & _T_7661; // @[lib.scala 393:57]
  wire  _T_7673 = _T_4970 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7674 = perr_ic_index_ff == 7'h46; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7676 = _T_7674 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7677 = _T_7673 | _T_7676; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7678 = _T_7677 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7681 = tag_valid_clken_2[0] & _T_7678; // @[lib.scala 393:57]
  wire  _T_7690 = _T_4971 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7691 = perr_ic_index_ff == 7'h47; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7693 = _T_7691 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7694 = _T_7690 | _T_7693; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7695 = _T_7694 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7698 = tag_valid_clken_2[0] & _T_7695; // @[lib.scala 393:57]
  wire  _T_7707 = _T_4972 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7708 = perr_ic_index_ff == 7'h48; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7710 = _T_7708 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7711 = _T_7707 | _T_7710; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7712 = _T_7711 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7715 = tag_valid_clken_2[0] & _T_7712; // @[lib.scala 393:57]
  wire  _T_7724 = _T_4973 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7725 = perr_ic_index_ff == 7'h49; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7727 = _T_7725 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7728 = _T_7724 | _T_7727; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7729 = _T_7728 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7732 = tag_valid_clken_2[0] & _T_7729; // @[lib.scala 393:57]
  wire  _T_7741 = _T_4974 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7742 = perr_ic_index_ff == 7'h4a; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7744 = _T_7742 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7745 = _T_7741 | _T_7744; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7746 = _T_7745 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7749 = tag_valid_clken_2[0] & _T_7746; // @[lib.scala 393:57]
  wire  _T_7758 = _T_4975 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7759 = perr_ic_index_ff == 7'h4b; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7761 = _T_7759 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7762 = _T_7758 | _T_7761; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7763 = _T_7762 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7766 = tag_valid_clken_2[0] & _T_7763; // @[lib.scala 393:57]
  wire  _T_7775 = _T_4976 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7776 = perr_ic_index_ff == 7'h4c; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7778 = _T_7776 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7779 = _T_7775 | _T_7778; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7780 = _T_7779 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7783 = tag_valid_clken_2[0] & _T_7780; // @[lib.scala 393:57]
  wire  _T_7792 = _T_4977 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7793 = perr_ic_index_ff == 7'h4d; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7795 = _T_7793 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7796 = _T_7792 | _T_7795; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7797 = _T_7796 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7800 = tag_valid_clken_2[0] & _T_7797; // @[lib.scala 393:57]
  wire  _T_7809 = _T_4978 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7810 = perr_ic_index_ff == 7'h4e; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7812 = _T_7810 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7813 = _T_7809 | _T_7812; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7814 = _T_7813 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7817 = tag_valid_clken_2[0] & _T_7814; // @[lib.scala 393:57]
  wire  _T_7826 = _T_4979 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7827 = perr_ic_index_ff == 7'h4f; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7829 = _T_7827 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7830 = _T_7826 | _T_7829; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7831 = _T_7830 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7834 = tag_valid_clken_2[0] & _T_7831; // @[lib.scala 393:57]
  wire  _T_7843 = _T_4980 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7844 = perr_ic_index_ff == 7'h50; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7846 = _T_7844 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7847 = _T_7843 | _T_7846; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7848 = _T_7847 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7851 = tag_valid_clken_2[0] & _T_7848; // @[lib.scala 393:57]
  wire  _T_7860 = _T_4981 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7861 = perr_ic_index_ff == 7'h51; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7863 = _T_7861 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7864 = _T_7860 | _T_7863; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7865 = _T_7864 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7868 = tag_valid_clken_2[0] & _T_7865; // @[lib.scala 393:57]
  wire  _T_7877 = _T_4982 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7878 = perr_ic_index_ff == 7'h52; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7880 = _T_7878 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7881 = _T_7877 | _T_7880; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7882 = _T_7881 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7885 = tag_valid_clken_2[0] & _T_7882; // @[lib.scala 393:57]
  wire  _T_7894 = _T_4983 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7895 = perr_ic_index_ff == 7'h53; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7897 = _T_7895 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7898 = _T_7894 | _T_7897; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7899 = _T_7898 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7902 = tag_valid_clken_2[0] & _T_7899; // @[lib.scala 393:57]
  wire  _T_7911 = _T_4984 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7912 = perr_ic_index_ff == 7'h54; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7914 = _T_7912 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7915 = _T_7911 | _T_7914; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7916 = _T_7915 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7919 = tag_valid_clken_2[0] & _T_7916; // @[lib.scala 393:57]
  wire  _T_7928 = _T_4985 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7929 = perr_ic_index_ff == 7'h55; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7931 = _T_7929 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7932 = _T_7928 | _T_7931; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7933 = _T_7932 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7936 = tag_valid_clken_2[0] & _T_7933; // @[lib.scala 393:57]
  wire  _T_7945 = _T_4986 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7946 = perr_ic_index_ff == 7'h56; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7948 = _T_7946 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7949 = _T_7945 | _T_7948; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7950 = _T_7949 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7953 = tag_valid_clken_2[0] & _T_7950; // @[lib.scala 393:57]
  wire  _T_7962 = _T_4987 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7963 = perr_ic_index_ff == 7'h57; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7965 = _T_7963 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7966 = _T_7962 | _T_7965; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7967 = _T_7966 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7970 = tag_valid_clken_2[0] & _T_7967; // @[lib.scala 393:57]
  wire  _T_7979 = _T_4988 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7980 = perr_ic_index_ff == 7'h58; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7982 = _T_7980 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_7983 = _T_7979 | _T_7982; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_7984 = _T_7983 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_7987 = tag_valid_clken_2[0] & _T_7984; // @[lib.scala 393:57]
  wire  _T_7996 = _T_4989 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_7997 = perr_ic_index_ff == 7'h59; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_7999 = _T_7997 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8000 = _T_7996 | _T_7999; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8001 = _T_8000 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8004 = tag_valid_clken_2[0] & _T_8001; // @[lib.scala 393:57]
  wire  _T_8013 = _T_4990 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8014 = perr_ic_index_ff == 7'h5a; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8016 = _T_8014 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8017 = _T_8013 | _T_8016; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8018 = _T_8017 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8021 = tag_valid_clken_2[0] & _T_8018; // @[lib.scala 393:57]
  wire  _T_8030 = _T_4991 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8031 = perr_ic_index_ff == 7'h5b; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8033 = _T_8031 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8034 = _T_8030 | _T_8033; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8035 = _T_8034 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8038 = tag_valid_clken_2[0] & _T_8035; // @[lib.scala 393:57]
  wire  _T_8047 = _T_4992 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8048 = perr_ic_index_ff == 7'h5c; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8050 = _T_8048 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8051 = _T_8047 | _T_8050; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8052 = _T_8051 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8055 = tag_valid_clken_2[0] & _T_8052; // @[lib.scala 393:57]
  wire  _T_8064 = _T_4993 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8065 = perr_ic_index_ff == 7'h5d; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8067 = _T_8065 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8068 = _T_8064 | _T_8067; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8069 = _T_8068 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8072 = tag_valid_clken_2[0] & _T_8069; // @[lib.scala 393:57]
  wire  _T_8081 = _T_4994 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8082 = perr_ic_index_ff == 7'h5e; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8084 = _T_8082 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8085 = _T_8081 | _T_8084; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8086 = _T_8085 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8089 = tag_valid_clken_2[0] & _T_8086; // @[lib.scala 393:57]
  wire  _T_8098 = _T_4995 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8099 = perr_ic_index_ff == 7'h5f; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8101 = _T_8099 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8102 = _T_8098 | _T_8101; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8103 = _T_8102 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8106 = tag_valid_clken_2[0] & _T_8103; // @[lib.scala 393:57]
  wire  _T_8115 = _T_4964 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8118 = _T_7572 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8119 = _T_8115 | _T_8118; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8120 = _T_8119 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8123 = tag_valid_clken_2[1] & _T_8120; // @[lib.scala 393:57]
  wire  _T_8132 = _T_4965 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8135 = _T_7589 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8136 = _T_8132 | _T_8135; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8137 = _T_8136 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8140 = tag_valid_clken_2[1] & _T_8137; // @[lib.scala 393:57]
  wire  _T_8149 = _T_4966 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8152 = _T_7606 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8153 = _T_8149 | _T_8152; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8154 = _T_8153 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8157 = tag_valid_clken_2[1] & _T_8154; // @[lib.scala 393:57]
  wire  _T_8166 = _T_4967 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8169 = _T_7623 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8170 = _T_8166 | _T_8169; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8171 = _T_8170 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8174 = tag_valid_clken_2[1] & _T_8171; // @[lib.scala 393:57]
  wire  _T_8183 = _T_4968 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8186 = _T_7640 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8187 = _T_8183 | _T_8186; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8188 = _T_8187 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8191 = tag_valid_clken_2[1] & _T_8188; // @[lib.scala 393:57]
  wire  _T_8200 = _T_4969 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8203 = _T_7657 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8204 = _T_8200 | _T_8203; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8205 = _T_8204 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8208 = tag_valid_clken_2[1] & _T_8205; // @[lib.scala 393:57]
  wire  _T_8217 = _T_4970 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8220 = _T_7674 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8221 = _T_8217 | _T_8220; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8222 = _T_8221 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8225 = tag_valid_clken_2[1] & _T_8222; // @[lib.scala 393:57]
  wire  _T_8234 = _T_4971 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8237 = _T_7691 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8238 = _T_8234 | _T_8237; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8239 = _T_8238 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8242 = tag_valid_clken_2[1] & _T_8239; // @[lib.scala 393:57]
  wire  _T_8251 = _T_4972 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8254 = _T_7708 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8255 = _T_8251 | _T_8254; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8256 = _T_8255 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8259 = tag_valid_clken_2[1] & _T_8256; // @[lib.scala 393:57]
  wire  _T_8268 = _T_4973 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8271 = _T_7725 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8272 = _T_8268 | _T_8271; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8273 = _T_8272 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8276 = tag_valid_clken_2[1] & _T_8273; // @[lib.scala 393:57]
  wire  _T_8285 = _T_4974 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8288 = _T_7742 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8289 = _T_8285 | _T_8288; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8290 = _T_8289 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8293 = tag_valid_clken_2[1] & _T_8290; // @[lib.scala 393:57]
  wire  _T_8302 = _T_4975 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8305 = _T_7759 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8306 = _T_8302 | _T_8305; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8307 = _T_8306 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8310 = tag_valid_clken_2[1] & _T_8307; // @[lib.scala 393:57]
  wire  _T_8319 = _T_4976 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8322 = _T_7776 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8323 = _T_8319 | _T_8322; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8324 = _T_8323 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8327 = tag_valid_clken_2[1] & _T_8324; // @[lib.scala 393:57]
  wire  _T_8336 = _T_4977 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8339 = _T_7793 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8340 = _T_8336 | _T_8339; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8341 = _T_8340 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8344 = tag_valid_clken_2[1] & _T_8341; // @[lib.scala 393:57]
  wire  _T_8353 = _T_4978 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8356 = _T_7810 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8357 = _T_8353 | _T_8356; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8358 = _T_8357 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8361 = tag_valid_clken_2[1] & _T_8358; // @[lib.scala 393:57]
  wire  _T_8370 = _T_4979 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8373 = _T_7827 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8374 = _T_8370 | _T_8373; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8375 = _T_8374 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8378 = tag_valid_clken_2[1] & _T_8375; // @[lib.scala 393:57]
  wire  _T_8387 = _T_4980 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8390 = _T_7844 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8391 = _T_8387 | _T_8390; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8392 = _T_8391 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8395 = tag_valid_clken_2[1] & _T_8392; // @[lib.scala 393:57]
  wire  _T_8404 = _T_4981 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8407 = _T_7861 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8408 = _T_8404 | _T_8407; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8409 = _T_8408 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8412 = tag_valid_clken_2[1] & _T_8409; // @[lib.scala 393:57]
  wire  _T_8421 = _T_4982 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8424 = _T_7878 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8425 = _T_8421 | _T_8424; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8426 = _T_8425 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8429 = tag_valid_clken_2[1] & _T_8426; // @[lib.scala 393:57]
  wire  _T_8438 = _T_4983 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8441 = _T_7895 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8442 = _T_8438 | _T_8441; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8443 = _T_8442 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8446 = tag_valid_clken_2[1] & _T_8443; // @[lib.scala 393:57]
  wire  _T_8455 = _T_4984 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8458 = _T_7912 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8459 = _T_8455 | _T_8458; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8460 = _T_8459 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8463 = tag_valid_clken_2[1] & _T_8460; // @[lib.scala 393:57]
  wire  _T_8472 = _T_4985 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8475 = _T_7929 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8476 = _T_8472 | _T_8475; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8477 = _T_8476 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8480 = tag_valid_clken_2[1] & _T_8477; // @[lib.scala 393:57]
  wire  _T_8489 = _T_4986 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8492 = _T_7946 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8493 = _T_8489 | _T_8492; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8494 = _T_8493 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8497 = tag_valid_clken_2[1] & _T_8494; // @[lib.scala 393:57]
  wire  _T_8506 = _T_4987 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8509 = _T_7963 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8510 = _T_8506 | _T_8509; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8511 = _T_8510 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8514 = tag_valid_clken_2[1] & _T_8511; // @[lib.scala 393:57]
  wire  _T_8523 = _T_4988 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8526 = _T_7980 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8527 = _T_8523 | _T_8526; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8528 = _T_8527 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8531 = tag_valid_clken_2[1] & _T_8528; // @[lib.scala 393:57]
  wire  _T_8540 = _T_4989 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8543 = _T_7997 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8544 = _T_8540 | _T_8543; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8545 = _T_8544 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8548 = tag_valid_clken_2[1] & _T_8545; // @[lib.scala 393:57]
  wire  _T_8557 = _T_4990 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8560 = _T_8014 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8561 = _T_8557 | _T_8560; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8562 = _T_8561 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8565 = tag_valid_clken_2[1] & _T_8562; // @[lib.scala 393:57]
  wire  _T_8574 = _T_4991 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8577 = _T_8031 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8578 = _T_8574 | _T_8577; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8579 = _T_8578 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8582 = tag_valid_clken_2[1] & _T_8579; // @[lib.scala 393:57]
  wire  _T_8591 = _T_4992 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8594 = _T_8048 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8595 = _T_8591 | _T_8594; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8596 = _T_8595 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8599 = tag_valid_clken_2[1] & _T_8596; // @[lib.scala 393:57]
  wire  _T_8608 = _T_4993 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8611 = _T_8065 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8612 = _T_8608 | _T_8611; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8613 = _T_8612 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8616 = tag_valid_clken_2[1] & _T_8613; // @[lib.scala 393:57]
  wire  _T_8625 = _T_4994 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8628 = _T_8082 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8629 = _T_8625 | _T_8628; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8630 = _T_8629 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8633 = tag_valid_clken_2[1] & _T_8630; // @[lib.scala 393:57]
  wire  _T_8642 = _T_4995 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8645 = _T_8099 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8646 = _T_8642 | _T_8645; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8647 = _T_8646 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8650 = tag_valid_clken_2[1] & _T_8647; // @[lib.scala 393:57]
  wire  _T_8659 = _T_4996 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8660 = perr_ic_index_ff == 7'h60; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8662 = _T_8660 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8663 = _T_8659 | _T_8662; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8664 = _T_8663 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8667 = tag_valid_clken_3[0] & _T_8664; // @[lib.scala 393:57]
  wire  _T_8676 = _T_4997 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8677 = perr_ic_index_ff == 7'h61; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8679 = _T_8677 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8680 = _T_8676 | _T_8679; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8681 = _T_8680 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8684 = tag_valid_clken_3[0] & _T_8681; // @[lib.scala 393:57]
  wire  _T_8693 = _T_4998 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8694 = perr_ic_index_ff == 7'h62; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8696 = _T_8694 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8697 = _T_8693 | _T_8696; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8698 = _T_8697 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8701 = tag_valid_clken_3[0] & _T_8698; // @[lib.scala 393:57]
  wire  _T_8710 = _T_4999 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8711 = perr_ic_index_ff == 7'h63; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8713 = _T_8711 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8714 = _T_8710 | _T_8713; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8715 = _T_8714 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8718 = tag_valid_clken_3[0] & _T_8715; // @[lib.scala 393:57]
  wire  _T_8727 = _T_5000 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8728 = perr_ic_index_ff == 7'h64; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8730 = _T_8728 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8731 = _T_8727 | _T_8730; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8732 = _T_8731 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8735 = tag_valid_clken_3[0] & _T_8732; // @[lib.scala 393:57]
  wire  _T_8744 = _T_5001 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8745 = perr_ic_index_ff == 7'h65; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8747 = _T_8745 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8748 = _T_8744 | _T_8747; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8749 = _T_8748 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8752 = tag_valid_clken_3[0] & _T_8749; // @[lib.scala 393:57]
  wire  _T_8761 = _T_5002 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8762 = perr_ic_index_ff == 7'h66; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8764 = _T_8762 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8765 = _T_8761 | _T_8764; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8766 = _T_8765 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8769 = tag_valid_clken_3[0] & _T_8766; // @[lib.scala 393:57]
  wire  _T_8778 = _T_5003 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8779 = perr_ic_index_ff == 7'h67; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8781 = _T_8779 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8782 = _T_8778 | _T_8781; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8783 = _T_8782 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8786 = tag_valid_clken_3[0] & _T_8783; // @[lib.scala 393:57]
  wire  _T_8795 = _T_5004 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8796 = perr_ic_index_ff == 7'h68; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8798 = _T_8796 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8799 = _T_8795 | _T_8798; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8800 = _T_8799 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8803 = tag_valid_clken_3[0] & _T_8800; // @[lib.scala 393:57]
  wire  _T_8812 = _T_5005 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8813 = perr_ic_index_ff == 7'h69; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8815 = _T_8813 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8816 = _T_8812 | _T_8815; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8817 = _T_8816 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8820 = tag_valid_clken_3[0] & _T_8817; // @[lib.scala 393:57]
  wire  _T_8829 = _T_5006 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8830 = perr_ic_index_ff == 7'h6a; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8832 = _T_8830 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8833 = _T_8829 | _T_8832; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8834 = _T_8833 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8837 = tag_valid_clken_3[0] & _T_8834; // @[lib.scala 393:57]
  wire  _T_8846 = _T_5007 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8847 = perr_ic_index_ff == 7'h6b; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8849 = _T_8847 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8850 = _T_8846 | _T_8849; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8851 = _T_8850 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8854 = tag_valid_clken_3[0] & _T_8851; // @[lib.scala 393:57]
  wire  _T_8863 = _T_5008 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8864 = perr_ic_index_ff == 7'h6c; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8866 = _T_8864 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8867 = _T_8863 | _T_8866; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8868 = _T_8867 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8871 = tag_valid_clken_3[0] & _T_8868; // @[lib.scala 393:57]
  wire  _T_8880 = _T_5009 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8881 = perr_ic_index_ff == 7'h6d; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8883 = _T_8881 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8884 = _T_8880 | _T_8883; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8885 = _T_8884 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8888 = tag_valid_clken_3[0] & _T_8885; // @[lib.scala 393:57]
  wire  _T_8897 = _T_5010 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8898 = perr_ic_index_ff == 7'h6e; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8900 = _T_8898 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8901 = _T_8897 | _T_8900; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8902 = _T_8901 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8905 = tag_valid_clken_3[0] & _T_8902; // @[lib.scala 393:57]
  wire  _T_8914 = _T_5011 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8915 = perr_ic_index_ff == 7'h6f; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8917 = _T_8915 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8918 = _T_8914 | _T_8917; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8919 = _T_8918 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8922 = tag_valid_clken_3[0] & _T_8919; // @[lib.scala 393:57]
  wire  _T_8931 = _T_5012 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8932 = perr_ic_index_ff == 7'h70; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8934 = _T_8932 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8935 = _T_8931 | _T_8934; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8936 = _T_8935 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8939 = tag_valid_clken_3[0] & _T_8936; // @[lib.scala 393:57]
  wire  _T_8948 = _T_5013 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8949 = perr_ic_index_ff == 7'h71; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8951 = _T_8949 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8952 = _T_8948 | _T_8951; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8953 = _T_8952 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8956 = tag_valid_clken_3[0] & _T_8953; // @[lib.scala 393:57]
  wire  _T_8965 = _T_5014 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8966 = perr_ic_index_ff == 7'h72; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8968 = _T_8966 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8969 = _T_8965 | _T_8968; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8970 = _T_8969 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8973 = tag_valid_clken_3[0] & _T_8970; // @[lib.scala 393:57]
  wire  _T_8982 = _T_5015 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_8983 = perr_ic_index_ff == 7'h73; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_8985 = _T_8983 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_8986 = _T_8982 | _T_8985; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_8987 = _T_8986 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_8990 = tag_valid_clken_3[0] & _T_8987; // @[lib.scala 393:57]
  wire  _T_8999 = _T_5016 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9000 = perr_ic_index_ff == 7'h74; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9002 = _T_9000 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9003 = _T_8999 | _T_9002; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9004 = _T_9003 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9007 = tag_valid_clken_3[0] & _T_9004; // @[lib.scala 393:57]
  wire  _T_9016 = _T_5017 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9017 = perr_ic_index_ff == 7'h75; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9019 = _T_9017 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9020 = _T_9016 | _T_9019; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9021 = _T_9020 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9024 = tag_valid_clken_3[0] & _T_9021; // @[lib.scala 393:57]
  wire  _T_9033 = _T_5018 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9034 = perr_ic_index_ff == 7'h76; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9036 = _T_9034 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9037 = _T_9033 | _T_9036; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9038 = _T_9037 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9041 = tag_valid_clken_3[0] & _T_9038; // @[lib.scala 393:57]
  wire  _T_9050 = _T_5019 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9051 = perr_ic_index_ff == 7'h77; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9053 = _T_9051 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9054 = _T_9050 | _T_9053; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9055 = _T_9054 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9058 = tag_valid_clken_3[0] & _T_9055; // @[lib.scala 393:57]
  wire  _T_9067 = _T_5020 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9068 = perr_ic_index_ff == 7'h78; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9070 = _T_9068 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9071 = _T_9067 | _T_9070; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9072 = _T_9071 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9075 = tag_valid_clken_3[0] & _T_9072; // @[lib.scala 393:57]
  wire  _T_9084 = _T_5021 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9085 = perr_ic_index_ff == 7'h79; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9087 = _T_9085 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9088 = _T_9084 | _T_9087; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9089 = _T_9088 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9092 = tag_valid_clken_3[0] & _T_9089; // @[lib.scala 393:57]
  wire  _T_9101 = _T_5022 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9102 = perr_ic_index_ff == 7'h7a; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9104 = _T_9102 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9105 = _T_9101 | _T_9104; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9106 = _T_9105 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9109 = tag_valid_clken_3[0] & _T_9106; // @[lib.scala 393:57]
  wire  _T_9118 = _T_5023 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9119 = perr_ic_index_ff == 7'h7b; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9121 = _T_9119 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9122 = _T_9118 | _T_9121; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9123 = _T_9122 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9126 = tag_valid_clken_3[0] & _T_9123; // @[lib.scala 393:57]
  wire  _T_9135 = _T_5024 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9136 = perr_ic_index_ff == 7'h7c; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9138 = _T_9136 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9139 = _T_9135 | _T_9138; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9140 = _T_9139 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9143 = tag_valid_clken_3[0] & _T_9140; // @[lib.scala 393:57]
  wire  _T_9152 = _T_5025 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9153 = perr_ic_index_ff == 7'h7d; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9155 = _T_9153 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9156 = _T_9152 | _T_9155; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9157 = _T_9156 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9160 = tag_valid_clken_3[0] & _T_9157; // @[lib.scala 393:57]
  wire  _T_9169 = _T_5026 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9170 = perr_ic_index_ff == 7'h7e; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9172 = _T_9170 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9173 = _T_9169 | _T_9172; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9174 = _T_9173 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9177 = tag_valid_clken_3[0] & _T_9174; // @[lib.scala 393:57]
  wire  _T_9186 = _T_5027 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9187 = perr_ic_index_ff == 7'h7f; // @[ifu_mem_ctl.scala 654:204]
  wire  _T_9189 = _T_9187 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9190 = _T_9186 | _T_9189; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9191 = _T_9190 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9194 = tag_valid_clken_3[0] & _T_9191; // @[lib.scala 393:57]
  wire  _T_9203 = _T_4996 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9206 = _T_8660 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9207 = _T_9203 | _T_9206; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9208 = _T_9207 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9211 = tag_valid_clken_3[1] & _T_9208; // @[lib.scala 393:57]
  wire  _T_9220 = _T_4997 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9223 = _T_8677 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9224 = _T_9220 | _T_9223; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9225 = _T_9224 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9228 = tag_valid_clken_3[1] & _T_9225; // @[lib.scala 393:57]
  wire  _T_9237 = _T_4998 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9240 = _T_8694 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9241 = _T_9237 | _T_9240; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9242 = _T_9241 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9245 = tag_valid_clken_3[1] & _T_9242; // @[lib.scala 393:57]
  wire  _T_9254 = _T_4999 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9257 = _T_8711 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9258 = _T_9254 | _T_9257; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9259 = _T_9258 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9262 = tag_valid_clken_3[1] & _T_9259; // @[lib.scala 393:57]
  wire  _T_9271 = _T_5000 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9274 = _T_8728 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9275 = _T_9271 | _T_9274; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9276 = _T_9275 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9279 = tag_valid_clken_3[1] & _T_9276; // @[lib.scala 393:57]
  wire  _T_9288 = _T_5001 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9291 = _T_8745 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9292 = _T_9288 | _T_9291; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9293 = _T_9292 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9296 = tag_valid_clken_3[1] & _T_9293; // @[lib.scala 393:57]
  wire  _T_9305 = _T_5002 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9308 = _T_8762 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9309 = _T_9305 | _T_9308; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9310 = _T_9309 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9313 = tag_valid_clken_3[1] & _T_9310; // @[lib.scala 393:57]
  wire  _T_9322 = _T_5003 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9325 = _T_8779 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9326 = _T_9322 | _T_9325; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9327 = _T_9326 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9330 = tag_valid_clken_3[1] & _T_9327; // @[lib.scala 393:57]
  wire  _T_9339 = _T_5004 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9342 = _T_8796 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9343 = _T_9339 | _T_9342; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9344 = _T_9343 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9347 = tag_valid_clken_3[1] & _T_9344; // @[lib.scala 393:57]
  wire  _T_9356 = _T_5005 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9359 = _T_8813 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9360 = _T_9356 | _T_9359; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9361 = _T_9360 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9364 = tag_valid_clken_3[1] & _T_9361; // @[lib.scala 393:57]
  wire  _T_9373 = _T_5006 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9376 = _T_8830 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9377 = _T_9373 | _T_9376; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9378 = _T_9377 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9381 = tag_valid_clken_3[1] & _T_9378; // @[lib.scala 393:57]
  wire  _T_9390 = _T_5007 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9393 = _T_8847 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9394 = _T_9390 | _T_9393; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9395 = _T_9394 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9398 = tag_valid_clken_3[1] & _T_9395; // @[lib.scala 393:57]
  wire  _T_9407 = _T_5008 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9410 = _T_8864 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9411 = _T_9407 | _T_9410; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9412 = _T_9411 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9415 = tag_valid_clken_3[1] & _T_9412; // @[lib.scala 393:57]
  wire  _T_9424 = _T_5009 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9427 = _T_8881 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9428 = _T_9424 | _T_9427; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9429 = _T_9428 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9432 = tag_valid_clken_3[1] & _T_9429; // @[lib.scala 393:57]
  wire  _T_9441 = _T_5010 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9444 = _T_8898 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9445 = _T_9441 | _T_9444; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9446 = _T_9445 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9449 = tag_valid_clken_3[1] & _T_9446; // @[lib.scala 393:57]
  wire  _T_9458 = _T_5011 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9461 = _T_8915 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9462 = _T_9458 | _T_9461; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9463 = _T_9462 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9466 = tag_valid_clken_3[1] & _T_9463; // @[lib.scala 393:57]
  wire  _T_9475 = _T_5012 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9478 = _T_8932 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9479 = _T_9475 | _T_9478; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9480 = _T_9479 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9483 = tag_valid_clken_3[1] & _T_9480; // @[lib.scala 393:57]
  wire  _T_9492 = _T_5013 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9495 = _T_8949 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9496 = _T_9492 | _T_9495; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9497 = _T_9496 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9500 = tag_valid_clken_3[1] & _T_9497; // @[lib.scala 393:57]
  wire  _T_9509 = _T_5014 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9512 = _T_8966 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9513 = _T_9509 | _T_9512; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9514 = _T_9513 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9517 = tag_valid_clken_3[1] & _T_9514; // @[lib.scala 393:57]
  wire  _T_9526 = _T_5015 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9529 = _T_8983 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9530 = _T_9526 | _T_9529; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9531 = _T_9530 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9534 = tag_valid_clken_3[1] & _T_9531; // @[lib.scala 393:57]
  wire  _T_9543 = _T_5016 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9546 = _T_9000 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9547 = _T_9543 | _T_9546; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9548 = _T_9547 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9551 = tag_valid_clken_3[1] & _T_9548; // @[lib.scala 393:57]
  wire  _T_9560 = _T_5017 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9563 = _T_9017 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9564 = _T_9560 | _T_9563; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9565 = _T_9564 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9568 = tag_valid_clken_3[1] & _T_9565; // @[lib.scala 393:57]
  wire  _T_9577 = _T_5018 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9580 = _T_9034 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9581 = _T_9577 | _T_9580; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9582 = _T_9581 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9585 = tag_valid_clken_3[1] & _T_9582; // @[lib.scala 393:57]
  wire  _T_9594 = _T_5019 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9597 = _T_9051 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9598 = _T_9594 | _T_9597; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9599 = _T_9598 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9602 = tag_valid_clken_3[1] & _T_9599; // @[lib.scala 393:57]
  wire  _T_9611 = _T_5020 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9614 = _T_9068 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9615 = _T_9611 | _T_9614; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9616 = _T_9615 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9619 = tag_valid_clken_3[1] & _T_9616; // @[lib.scala 393:57]
  wire  _T_9628 = _T_5021 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9631 = _T_9085 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9632 = _T_9628 | _T_9631; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9633 = _T_9632 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9636 = tag_valid_clken_3[1] & _T_9633; // @[lib.scala 393:57]
  wire  _T_9645 = _T_5022 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9648 = _T_9102 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9649 = _T_9645 | _T_9648; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9650 = _T_9649 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9653 = tag_valid_clken_3[1] & _T_9650; // @[lib.scala 393:57]
  wire  _T_9662 = _T_5023 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9665 = _T_9119 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9666 = _T_9662 | _T_9665; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9667 = _T_9666 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9670 = tag_valid_clken_3[1] & _T_9667; // @[lib.scala 393:57]
  wire  _T_9679 = _T_5024 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9682 = _T_9136 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9683 = _T_9679 | _T_9682; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9684 = _T_9683 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9687 = tag_valid_clken_3[1] & _T_9684; // @[lib.scala 393:57]
  wire  _T_9696 = _T_5025 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9699 = _T_9153 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9700 = _T_9696 | _T_9699; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9701 = _T_9700 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9704 = tag_valid_clken_3[1] & _T_9701; // @[lib.scala 393:57]
  wire  _T_9713 = _T_5026 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9716 = _T_9170 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9717 = _T_9713 | _T_9716; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9718 = _T_9717 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9721 = tag_valid_clken_3[1] & _T_9718; // @[lib.scala 393:57]
  wire  _T_9730 = _T_5027 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 654:161]
  wire  _T_9733 = _T_9187 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 654:226]
  wire  _T_9734 = _T_9730 | _T_9733; // @[ifu_mem_ctl.scala 654:183]
  wire  _T_9735 = _T_9734 | reset_all_tags; // @[ifu_mem_ctl.scala 654:249]
  wire  _T_9738 = tag_valid_clken_3[1] & _T_9735; // @[lib.scala 393:57]
  wire  _T_10539 = ~fetch_uncacheable_ff; // @[ifu_mem_ctl.scala 702:63]
  wire  _T_10540 = _T_10539 & ifc_fetch_req_f_raw; // @[ifu_mem_ctl.scala 702:85]
  wire [1:0] _T_10542 = _T_10540 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10552; // @[Reg.scala 27:20]
  wire  _T_10550 = ic_act_miss_f ^ _T_10552; // @[lib.scala 475:21]
  wire  _T_10551 = |_T_10550; // @[lib.scala 475:29]
  reg  _T_10556; // @[Reg.scala 27:20]
  wire  _T_10554 = ic_act_hit_f ^ _T_10556; // @[lib.scala 475:21]
  wire  _T_10555 = |_T_10554; // @[lib.scala 475:29]
  reg  _T_10561; // @[Reg.scala 27:20]
  wire  _T_10559 = _T_2500 ^ _T_10561; // @[lib.scala 475:21]
  wire  _T_10560 = |_T_10559; // @[lib.scala 475:29]
  wire  _T_10562 = ~ifu_bus_arready_ff; // @[ifu_mem_ctl.scala 710:69]
  wire  _T_10563 = ifu_bus_arvalid_ff & _T_10562; // @[ifu_mem_ctl.scala 710:67]
  wire  _T_10564 = _T_10563 & miss_pending; // @[ifu_mem_ctl.scala 710:89]
  reg  _T_10568; // @[Reg.scala 27:20]
  wire  _T_10566 = _T_10564 ^ _T_10568; // @[lib.scala 475:21]
  wire  _T_10567 = |_T_10566; // @[lib.scala 475:29]
  reg  _T_10572; // @[Reg.scala 27:20]
  wire  _T_10570 = bus_cmd_sent ^ _T_10572; // @[lib.scala 475:21]
  wire  _T_10571 = |_T_10570; // @[lib.scala 475:29]
  wire  _T_10575 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[ifu_mem_ctl.scala 718:84]
  wire  _T_10577 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[ifu_mem_ctl.scala 718:150]
  wire  _T_10579 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[ifu_mem_ctl.scala 719:63]
  wire  _T_10581 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[ifu_mem_ctl.scala 719:129]
  wire [3:0] _T_10584 = {_T_10575,_T_10577,_T_10579,_T_10581}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[ifu_mem_ctl.scala 721:53]
  wire  _T_10592 = io_ic_debug_rd_en ^ ic_debug_rd_en_ff; // @[lib.scala 475:21]
  wire  _T_10593 = |_T_10592; // @[lib.scala 475:29]
  reg  _T_10598; // @[Reg.scala 27:20]
  wire  _T_10596 = ic_debug_rd_en_ff ^ _T_10598; // @[lib.scala 475:21]
  wire  _T_10597 = |_T_10596; // @[lib.scala 475:29]
  wire  _T_10660 = ifc_region_acc_fault_memory_bf ^ ifc_region_acc_fault_memory_f; // @[lib.scala 475:21]
  wire  _T_10661 = |_T_10660; // @[lib.scala 475:29]
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en)
  );
  rvclkhdr rvclkhdr_20 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en)
  );
  rvclkhdr rvclkhdr_21 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en)
  );
  rvclkhdr rvclkhdr_22 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en)
  );
  rvclkhdr rvclkhdr_23 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en)
  );
  rvclkhdr rvclkhdr_24 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en)
  );
  rvclkhdr rvclkhdr_25 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en)
  );
  rvclkhdr rvclkhdr_26 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en)
  );
  rvclkhdr rvclkhdr_27 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en)
  );
  rvclkhdr rvclkhdr_28 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en)
  );
  rvclkhdr rvclkhdr_29 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en)
  );
  rvclkhdr rvclkhdr_30 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en)
  );
  rvclkhdr rvclkhdr_31 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en)
  );
  rvclkhdr rvclkhdr_32 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en)
  );
  rvclkhdr rvclkhdr_33 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en)
  );
  rvclkhdr rvclkhdr_34 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en)
  );
  rvclkhdr rvclkhdr_35 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en)
  );
  rvclkhdr rvclkhdr_36 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en)
  );
  rvclkhdr rvclkhdr_37 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en)
  );
  rvclkhdr rvclkhdr_38 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en)
  );
  rvclkhdr rvclkhdr_39 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en)
  );
  rvclkhdr rvclkhdr_40 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en)
  );
  rvclkhdr rvclkhdr_41 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en)
  );
  rvclkhdr rvclkhdr_42 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en)
  );
  rvclkhdr rvclkhdr_43 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en)
  );
  rvclkhdr rvclkhdr_44 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en)
  );
  rvclkhdr rvclkhdr_45 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en)
  );
  rvclkhdr rvclkhdr_46 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en)
  );
  assign io_dec_mem_ctrl_ifu_pmu_ic_miss = _T_10552; // @[ifu_mem_ctl.scala 707:37]
  assign io_dec_mem_ctrl_ifu_pmu_ic_hit = _T_10556; // @[ifu_mem_ctl.scala 708:37]
  assign io_dec_mem_ctrl_ifu_pmu_bus_error = _T_10561; // @[ifu_mem_ctl.scala 709:37]
  assign io_dec_mem_ctrl_ifu_pmu_bus_busy = _T_10568; // @[ifu_mem_ctl.scala 710:37]
  assign io_dec_mem_ctrl_ifu_pmu_bus_trxn = _T_10572; // @[ifu_mem_ctl.scala 711:37]
  assign io_dec_mem_ctrl_ifu_ic_error_start = _T_1225 | ic_rd_parity_final_err; // @[ifu_mem_ctl.scala 252:38]
  assign io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err = _T_3981 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 571:48]
  assign io_dec_mem_ctrl_ifu_ic_debug_rd_data = _T_1237; // @[ifu_mem_ctl.scala 260:40]
  assign io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid = _T_10598; // @[ifu_mem_ctl.scala 725:46]
  assign io_dec_mem_ctrl_ifu_miss_state_idle = miss_state == 3'h0; // @[ifu_mem_ctl.scala 232:39]
  assign io_ifu_axi_ar_valid = ifu_bus_cmd_valid; // @[ifu_mem_ctl.scala 468:14 ifu_mem_ctl.scala 470:23]
  assign io_ifu_axi_ar_bits_id = bus_rd_addr_count & _T_2639; // @[ifu_mem_ctl.scala 468:14 ifu_mem_ctl.scala 471:25]
  assign io_ifu_axi_ar_bits_addr = _T_2641 & _T_2643; // @[ifu_mem_ctl.scala 468:14 ifu_mem_ctl.scala 472:27]
  assign io_ifu_axi_ar_bits_region = ifu_ic_req_addr_f[28:25]; // @[ifu_mem_ctl.scala 468:14 ifu_mem_ctl.scala 475:29]
  assign io_ifu_axi_r_ready = 1'h1; // @[ifu_mem_ctl.scala 468:14 ifu_mem_ctl.scala 477:22]
  assign io_iccm_rw_addr = _T_3180 ? io_dma_mem_ctl_dma_mem_addr[15:1] : _T_3187; // @[ifu_mem_ctl.scala 558:19]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2519; // @[ifu_mem_ctl.scala 385:27]
  assign io_iccm_correction_state = _T_2547 ? 1'h0 : _GEN_81; // @[ifu_mem_ctl.scala 419:28 ifu_mem_ctl.scala 431:32 ifu_mem_ctl.scala 438:32 ifu_mem_ctl.scala 445:32]
  assign io_iccm_wren = _T_2760 | iccm_correct_ecc; // @[ifu_mem_ctl.scala 532:16]
  assign io_iccm_rden = _T_2764 | _T_2765; // @[ifu_mem_ctl.scala 533:16]
  assign io_iccm_wr_size = _T_2770 & io_dma_mem_ctl_dma_mem_sz; // @[ifu_mem_ctl.scala 535:19]
  assign io_iccm_wr_data = _T_3142 ? _T_3143 : _T_3150; // @[ifu_mem_ctl.scala 539:19]
  assign io_ic_rw_addr = _T_360 | _T_361; // @[ifu_mem_ctl.scala 236:17]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10542; // @[ifu_mem_ctl.scala 702:19]
  assign io_ic_wr_en = bus_ic_wr_en & _T_4063; // @[ifu_mem_ctl.scala 601:15]
  assign io_ic_rd_en = _T_4055 | _T_4060; // @[ifu_mem_ctl.scala 592:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[ifu_mem_ctl.scala 249:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[ifu_mem_ctl.scala 249:17]
  assign io_ic_debug_wr_data = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[ifu_mem_ctl.scala 250:23]
  assign io_ic_debug_addr = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[ifu_mem_ctl.scala 714:20]
  assign io_ic_debug_rd_en = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[ifu_mem_ctl.scala 716:21]
  assign io_ic_debug_wr_en = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[ifu_mem_ctl.scala 717:21]
  assign io_ic_debug_tag_array = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[ifu_mem_ctl.scala 715:25]
  assign io_ic_debug_way = _T_10584[1:0]; // @[ifu_mem_ctl.scala 718:19]
  assign io_ic_premux_data = ic_premux_data_temp[63:0]; // @[ifu_mem_ctl.scala 287:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | _T_1280; // @[ifu_mem_ctl.scala 288:25]
  assign io_ifu_ic_mb_empty = _T_348 | _T_237; // @[ifu_mem_ctl.scala 231:22]
  assign io_ic_dma_active = _T_14 | io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu_mem_ctl.scala 93:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_4077; // @[ifu_mem_ctl.scala 602:21]
  assign io_iccm_dma_ecc_error = iccm_dma_ecc_error; // @[ifu_mem_ctl.scala 554:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid_temp; // @[ifu_mem_ctl.scala 552:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata_temp; // @[ifu_mem_ctl.scala 556:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag_temp; // @[ifu_mem_ctl.scala 548:20]
  assign io_iccm_ready = _T_2752 & _T_2742; // @[ifu_mem_ctl.scala 530:18]
  assign io_iccm_rd_ecc_double_err = _T_2153 ? _T_3990 : _T_3996; // @[ifu_mem_ctl.scala 572:31]
  assign io_iccm_dma_sb_error = _T_6 & dma_iccm_req_f; // @[ifu_mem_ctl.scala 91:24]
  assign io_ic_hit_f = _T_269 | _T_270; // @[ifu_mem_ctl.scala 191:15]
  assign io_ic_access_fault_f = _T_1302 & _T_1305; // @[ifu_mem_ctl.scala 293:24]
  assign io_ic_access_fault_type_f = _T_1307 ? 2'h1 : _T_1310; // @[ifu_mem_ctl.scala 294:29]
  assign io_ifu_async_error_start = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err | io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu_mem_ctl.scala 92:28]
  assign io_ic_fetch_val_f = {_T_1318,fetch_req_f_qual}; // @[ifu_mem_ctl.scala 296:21]
  assign io_ic_data_f = ic_final_data[31:0]; // @[ifu_mem_ctl.scala 290:16]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = ic_debug_rd_en_ff; // @[lib.scala 345:16]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_1_io_en = io_ifu_bus_clk_en & io_ifu_axi_r_valid; // @[lib.scala 412:17]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_2_io_en = ic_debug_rd_en_ff; // @[lib.scala 412:17]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_3_io_en = bus_ifu_wr_en & _T_1321; // @[lib.scala 412:17]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_4_io_en = bus_ifu_wr_en & _T_1321; // @[lib.scala 412:17]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_5_io_en = bus_ifu_wr_en & _T_1322; // @[lib.scala 412:17]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_6_io_en = bus_ifu_wr_en & _T_1322; // @[lib.scala 412:17]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_7_io_en = bus_ifu_wr_en & _T_1323; // @[lib.scala 412:17]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_8_io_en = bus_ifu_wr_en & _T_1323; // @[lib.scala 412:17]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_9_io_en = bus_ifu_wr_en & _T_1324; // @[lib.scala 412:17]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_10_io_en = bus_ifu_wr_en & _T_1324; // @[lib.scala 412:17]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_11_io_en = bus_ifu_wr_en & _T_1325; // @[lib.scala 412:17]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_12_io_en = bus_ifu_wr_en & _T_1325; // @[lib.scala 412:17]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_13_io_en = bus_ifu_wr_en & _T_1326; // @[lib.scala 412:17]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_14_io_en = bus_ifu_wr_en & _T_1326; // @[lib.scala 412:17]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_15_io_en = bus_ifu_wr_en & _T_1327; // @[lib.scala 412:17]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_16_io_en = bus_ifu_wr_en & _T_1327; // @[lib.scala 412:17]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_17_io_en = bus_ifu_wr_en & _T_1328; // @[lib.scala 412:17]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_18_io_en = bus_ifu_wr_en & _T_1328; // @[lib.scala 412:17]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_19_io_en = _T_2521 & perr_state_en; // @[lib.scala 412:17]
  assign rvclkhdr_20_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_20_io_en = iccm_dma_rvalid_in; // @[lib.scala 412:17]
  assign rvclkhdr_21_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_21_io_en = _T_4008 | io_iccm_dma_sb_error; // @[lib.scala 412:17]
  assign rvclkhdr_22_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_22_io_en = _T_4008 | io_iccm_dma_sb_error; // @[lib.scala 412:17]
  assign rvclkhdr_23_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_23_io_en = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[lib.scala 345:16]
  assign rvclkhdr_24_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_24_io_en = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[lib.scala 345:16]
  assign rvclkhdr_25_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_25_io_en = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[lib.scala 345:16]
  assign rvclkhdr_26_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_26_io_en = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[lib.scala 345:16]
  assign rvclkhdr_27_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_27_io_en = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[lib.scala 345:16]
  assign rvclkhdr_28_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_28_io_en = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[lib.scala 345:16]
  assign rvclkhdr_29_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_29_io_en = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[lib.scala 345:16]
  assign rvclkhdr_30_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_30_io_en = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[lib.scala 345:16]
  assign rvclkhdr_31_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_31_io_en = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[lib.scala 345:16]
  assign rvclkhdr_32_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_32_io_en = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[lib.scala 345:16]
  assign rvclkhdr_33_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_33_io_en = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[lib.scala 345:16]
  assign rvclkhdr_34_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_34_io_en = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[lib.scala 345:16]
  assign rvclkhdr_35_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_35_io_en = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[lib.scala 345:16]
  assign rvclkhdr_36_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_36_io_en = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[lib.scala 345:16]
  assign rvclkhdr_37_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_37_io_en = ifu_status_wr_addr_ff[6:3] == 4'he; // @[lib.scala 345:16]
  assign rvclkhdr_38_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_38_io_en = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[lib.scala 345:16]
  assign rvclkhdr_39_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_39_io_en = tag_valid_clken_0[0]; // @[lib.scala 345:16]
  assign rvclkhdr_40_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_40_io_en = tag_valid_clken_0[1]; // @[lib.scala 345:16]
  assign rvclkhdr_41_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_41_io_en = tag_valid_clken_1[0]; // @[lib.scala 345:16]
  assign rvclkhdr_42_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_42_io_en = tag_valid_clken_1[1]; // @[lib.scala 345:16]
  assign rvclkhdr_43_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_43_io_en = tag_valid_clken_2[0]; // @[lib.scala 345:16]
  assign rvclkhdr_44_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_44_io_en = tag_valid_clken_2[1]; // @[lib.scala 345:16]
  assign rvclkhdr_45_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_45_io_en = tag_valid_clken_3[0]; // @[lib.scala 345:16]
  assign rvclkhdr_46_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_46_io_en = tag_valid_clken_3[1]; // @[lib.scala 345:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_11 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_17 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_18 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_19 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_20 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_21 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_23 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_24 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_25 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_26 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_27 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_29 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_30 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_32 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_33 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_34 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_35 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_36 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_37 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_38 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_39 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_40 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_41 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_42 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_43 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_44 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_45 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_46 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_47 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_48 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_49 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_50 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_51 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_52 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_53 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_54 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_55 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_56 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_57 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_58 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_59 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_60 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_61 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_62 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_63 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_64 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_65 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_66 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_67 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_68 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_69 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_70 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_71 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_72 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_73 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_74 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_75 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_76 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_77 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_78 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_79 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_80 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_81 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_82 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_83 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_84 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_85 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_86 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_87 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_88 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_89 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_90 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_91 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_92 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_93 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_94 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_95 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_96 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_97 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_98 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_99 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_100 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_101 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_102 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_103 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_104 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_105 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_106 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_107 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_108 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_109 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_110 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_111 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_112 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_113 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_114 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_115 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_116 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_117 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_118 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_119 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_120 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_121 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_out_122 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way_status_out_123 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way_status_out_124 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way_status_out_125 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way_status_out_126 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way_status_out_127 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagv_mb_scnd_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_152[30:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  reset_ic_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  miss_addr = _RAND_160[25:0];
  _RAND_161 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_441[0:0];
  _RAND_442 = {3{`RANDOM}};
  _T_1237 = _RAND_442[70:0];
  _RAND_443 = {1{`RANDOM}};
  ifc_region_acc_fault_memory_f = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_444[6:0];
  _RAND_445 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  bus_cmd_req_hold = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_448[2:0];
  _RAND_449 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_451[0:0];
  _RAND_452 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_452[38:0];
  _RAND_453 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_454[2:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_dma_rtag_temp = _RAND_455[2:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_dma_rvalid_temp = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_dma_ecc_error = _RAND_457[0:0];
  _RAND_458 = {2{`RANDOM}};
  iccm_dma_rdata_temp = _RAND_458[63:0];
  _RAND_459 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_459[13:0];
  _RAND_460 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_461[13:0];
  _RAND_462 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_462[6:0];
  _RAND_463 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  way_status_new_ff = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  ic_valid_ff = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_10552 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_10556 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_10561 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  _T_10568 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  _T_10572 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  _T_10598 = _RAND_472[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    flush_final_f = 1'h0;
  end
  if (reset) begin
    ifc_fetch_req_f_raw = 1'h0;
  end
  if (reset) begin
    miss_state = 3'h0;
  end
  if (reset) begin
    scnd_miss_req_q = 1'h0;
  end
  if (reset) begin
    ifu_fetch_addr_int_f = 31'h0;
  end
  if (reset) begin
    ifc_iccm_access_f = 1'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_in = 1'h0;
  end
  if (reset) begin
    dma_iccm_req_f = 1'h0;
  end
  if (reset) begin
    perr_state = 3'h0;
  end
  if (reset) begin
    err_stop_state = 2'h0;
  end
  if (reset) begin
    reset_all_tags = 1'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_final_f = 1'h0;
  end
  if (reset) begin
    ifu_bus_rvalid_unq_ff = 1'h0;
  end
  if (reset) begin
    bus_ifu_bus_clk_en_ff = 1'h0;
  end
  if (reset) begin
    uncacheable_miss_ff = 1'h0;
  end
  if (reset) begin
    bus_data_beat_count = 3'h0;
  end
  if (reset) begin
    ic_miss_buff_data_valid = 8'h0;
  end
  if (reset) begin
    imb_ff = 31'h0;
  end
  if (reset) begin
    last_data_recieved_ff = 1'h0;
  end
  if (reset) begin
    sel_mb_addr_ff = 1'h0;
  end
  if (reset) begin
    way_status_mb_scnd_ff = 1'h0;
  end
  if (reset) begin
    ifu_ic_rw_int_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_out_0 = 1'h0;
  end
  if (reset) begin
    way_status_out_1 = 1'h0;
  end
  if (reset) begin
    way_status_out_2 = 1'h0;
  end
  if (reset) begin
    way_status_out_3 = 1'h0;
  end
  if (reset) begin
    way_status_out_4 = 1'h0;
  end
  if (reset) begin
    way_status_out_5 = 1'h0;
  end
  if (reset) begin
    way_status_out_6 = 1'h0;
  end
  if (reset) begin
    way_status_out_7 = 1'h0;
  end
  if (reset) begin
    way_status_out_8 = 1'h0;
  end
  if (reset) begin
    way_status_out_9 = 1'h0;
  end
  if (reset) begin
    way_status_out_10 = 1'h0;
  end
  if (reset) begin
    way_status_out_11 = 1'h0;
  end
  if (reset) begin
    way_status_out_12 = 1'h0;
  end
  if (reset) begin
    way_status_out_13 = 1'h0;
  end
  if (reset) begin
    way_status_out_14 = 1'h0;
  end
  if (reset) begin
    way_status_out_15 = 1'h0;
  end
  if (reset) begin
    way_status_out_16 = 1'h0;
  end
  if (reset) begin
    way_status_out_17 = 1'h0;
  end
  if (reset) begin
    way_status_out_18 = 1'h0;
  end
  if (reset) begin
    way_status_out_19 = 1'h0;
  end
  if (reset) begin
    way_status_out_20 = 1'h0;
  end
  if (reset) begin
    way_status_out_21 = 1'h0;
  end
  if (reset) begin
    way_status_out_22 = 1'h0;
  end
  if (reset) begin
    way_status_out_23 = 1'h0;
  end
  if (reset) begin
    way_status_out_24 = 1'h0;
  end
  if (reset) begin
    way_status_out_25 = 1'h0;
  end
  if (reset) begin
    way_status_out_26 = 1'h0;
  end
  if (reset) begin
    way_status_out_27 = 1'h0;
  end
  if (reset) begin
    way_status_out_28 = 1'h0;
  end
  if (reset) begin
    way_status_out_29 = 1'h0;
  end
  if (reset) begin
    way_status_out_30 = 1'h0;
  end
  if (reset) begin
    way_status_out_31 = 1'h0;
  end
  if (reset) begin
    way_status_out_32 = 1'h0;
  end
  if (reset) begin
    way_status_out_33 = 1'h0;
  end
  if (reset) begin
    way_status_out_34 = 1'h0;
  end
  if (reset) begin
    way_status_out_35 = 1'h0;
  end
  if (reset) begin
    way_status_out_36 = 1'h0;
  end
  if (reset) begin
    way_status_out_37 = 1'h0;
  end
  if (reset) begin
    way_status_out_38 = 1'h0;
  end
  if (reset) begin
    way_status_out_39 = 1'h0;
  end
  if (reset) begin
    way_status_out_40 = 1'h0;
  end
  if (reset) begin
    way_status_out_41 = 1'h0;
  end
  if (reset) begin
    way_status_out_42 = 1'h0;
  end
  if (reset) begin
    way_status_out_43 = 1'h0;
  end
  if (reset) begin
    way_status_out_44 = 1'h0;
  end
  if (reset) begin
    way_status_out_45 = 1'h0;
  end
  if (reset) begin
    way_status_out_46 = 1'h0;
  end
  if (reset) begin
    way_status_out_47 = 1'h0;
  end
  if (reset) begin
    way_status_out_48 = 1'h0;
  end
  if (reset) begin
    way_status_out_49 = 1'h0;
  end
  if (reset) begin
    way_status_out_50 = 1'h0;
  end
  if (reset) begin
    way_status_out_51 = 1'h0;
  end
  if (reset) begin
    way_status_out_52 = 1'h0;
  end
  if (reset) begin
    way_status_out_53 = 1'h0;
  end
  if (reset) begin
    way_status_out_54 = 1'h0;
  end
  if (reset) begin
    way_status_out_55 = 1'h0;
  end
  if (reset) begin
    way_status_out_56 = 1'h0;
  end
  if (reset) begin
    way_status_out_57 = 1'h0;
  end
  if (reset) begin
    way_status_out_58 = 1'h0;
  end
  if (reset) begin
    way_status_out_59 = 1'h0;
  end
  if (reset) begin
    way_status_out_60 = 1'h0;
  end
  if (reset) begin
    way_status_out_61 = 1'h0;
  end
  if (reset) begin
    way_status_out_62 = 1'h0;
  end
  if (reset) begin
    way_status_out_63 = 1'h0;
  end
  if (reset) begin
    way_status_out_64 = 1'h0;
  end
  if (reset) begin
    way_status_out_65 = 1'h0;
  end
  if (reset) begin
    way_status_out_66 = 1'h0;
  end
  if (reset) begin
    way_status_out_67 = 1'h0;
  end
  if (reset) begin
    way_status_out_68 = 1'h0;
  end
  if (reset) begin
    way_status_out_69 = 1'h0;
  end
  if (reset) begin
    way_status_out_70 = 1'h0;
  end
  if (reset) begin
    way_status_out_71 = 1'h0;
  end
  if (reset) begin
    way_status_out_72 = 1'h0;
  end
  if (reset) begin
    way_status_out_73 = 1'h0;
  end
  if (reset) begin
    way_status_out_74 = 1'h0;
  end
  if (reset) begin
    way_status_out_75 = 1'h0;
  end
  if (reset) begin
    way_status_out_76 = 1'h0;
  end
  if (reset) begin
    way_status_out_77 = 1'h0;
  end
  if (reset) begin
    way_status_out_78 = 1'h0;
  end
  if (reset) begin
    way_status_out_79 = 1'h0;
  end
  if (reset) begin
    way_status_out_80 = 1'h0;
  end
  if (reset) begin
    way_status_out_81 = 1'h0;
  end
  if (reset) begin
    way_status_out_82 = 1'h0;
  end
  if (reset) begin
    way_status_out_83 = 1'h0;
  end
  if (reset) begin
    way_status_out_84 = 1'h0;
  end
  if (reset) begin
    way_status_out_85 = 1'h0;
  end
  if (reset) begin
    way_status_out_86 = 1'h0;
  end
  if (reset) begin
    way_status_out_87 = 1'h0;
  end
  if (reset) begin
    way_status_out_88 = 1'h0;
  end
  if (reset) begin
    way_status_out_89 = 1'h0;
  end
  if (reset) begin
    way_status_out_90 = 1'h0;
  end
  if (reset) begin
    way_status_out_91 = 1'h0;
  end
  if (reset) begin
    way_status_out_92 = 1'h0;
  end
  if (reset) begin
    way_status_out_93 = 1'h0;
  end
  if (reset) begin
    way_status_out_94 = 1'h0;
  end
  if (reset) begin
    way_status_out_95 = 1'h0;
  end
  if (reset) begin
    way_status_out_96 = 1'h0;
  end
  if (reset) begin
    way_status_out_97 = 1'h0;
  end
  if (reset) begin
    way_status_out_98 = 1'h0;
  end
  if (reset) begin
    way_status_out_99 = 1'h0;
  end
  if (reset) begin
    way_status_out_100 = 1'h0;
  end
  if (reset) begin
    way_status_out_101 = 1'h0;
  end
  if (reset) begin
    way_status_out_102 = 1'h0;
  end
  if (reset) begin
    way_status_out_103 = 1'h0;
  end
  if (reset) begin
    way_status_out_104 = 1'h0;
  end
  if (reset) begin
    way_status_out_105 = 1'h0;
  end
  if (reset) begin
    way_status_out_106 = 1'h0;
  end
  if (reset) begin
    way_status_out_107 = 1'h0;
  end
  if (reset) begin
    way_status_out_108 = 1'h0;
  end
  if (reset) begin
    way_status_out_109 = 1'h0;
  end
  if (reset) begin
    way_status_out_110 = 1'h0;
  end
  if (reset) begin
    way_status_out_111 = 1'h0;
  end
  if (reset) begin
    way_status_out_112 = 1'h0;
  end
  if (reset) begin
    way_status_out_113 = 1'h0;
  end
  if (reset) begin
    way_status_out_114 = 1'h0;
  end
  if (reset) begin
    way_status_out_115 = 1'h0;
  end
  if (reset) begin
    way_status_out_116 = 1'h0;
  end
  if (reset) begin
    way_status_out_117 = 1'h0;
  end
  if (reset) begin
    way_status_out_118 = 1'h0;
  end
  if (reset) begin
    way_status_out_119 = 1'h0;
  end
  if (reset) begin
    way_status_out_120 = 1'h0;
  end
  if (reset) begin
    way_status_out_121 = 1'h0;
  end
  if (reset) begin
    way_status_out_122 = 1'h0;
  end
  if (reset) begin
    way_status_out_123 = 1'h0;
  end
  if (reset) begin
    way_status_out_124 = 1'h0;
  end
  if (reset) begin
    way_status_out_125 = 1'h0;
  end
  if (reset) begin
    way_status_out_126 = 1'h0;
  end
  if (reset) begin
    way_status_out_127 = 1'h0;
  end
  if (reset) begin
    tagv_mb_scnd_ff = 2'h0;
  end
  if (reset) begin
    uncacheable_miss_scnd_ff = 1'h0;
  end
  if (reset) begin
    imb_scnd_ff = 31'h0;
  end
  if (reset) begin
    ifu_bus_rid_ff = 3'h0;
  end
  if (reset) begin
    ifu_bus_rresp_ff = 2'h0;
  end
  if (reset) begin
    ifu_wr_data_comb_err_ff = 1'h0;
  end
  if (reset) begin
    way_status_mb_ff = 1'h0;
  end
  if (reset) begin
    tagv_mb_ff = 2'h0;
  end
  if (reset) begin
    reset_ic_ff = 1'h0;
  end
  if (reset) begin
    fetch_uncacheable_ff = 1'h0;
  end
  if (reset) begin
    miss_addr = 26'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_f = 1'h0;
  end
  if (reset) begin
    bus_rd_addr_count = 3'h0;
  end
  if (reset) begin
    ic_act_miss_f_delayed = 1'h0;
  end
  if (reset) begin
    ifu_bus_rdata_ff = 64'h0;
  end
  if (reset) begin
    ic_miss_buff_data_0 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_1 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_2 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_3 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_4 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_5 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_6 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_7 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_8 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_9 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_10 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_11 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_12 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_13 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_14 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_15 = 32'h0;
  end
  if (reset) begin
    ic_crit_wd_rdy_new_ff = 1'h0;
  end
  if (reset) begin
    ic_miss_buff_data_error = 8'h0;
  end
  if (reset) begin
    ic_debug_ict_array_sel_ff = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_127 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_127 = 1'h0;
  end
  if (reset) begin
    ic_debug_way_ff = 2'h0;
  end
  if (reset) begin
    ic_debug_rd_en_ff = 1'h0;
  end
  if (reset) begin
    _T_1237 = 71'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_memory_f = 1'h0;
  end
  if (reset) begin
    perr_ic_index_ff = 7'h0;
  end
  if (reset) begin
    dma_sb_err_state_ff = 1'h0;
  end
  if (reset) begin
    bus_cmd_req_hold = 1'h0;
  end
  if (reset) begin
    ifu_bus_cmd_valid = 1'h0;
  end
  if (reset) begin
    bus_cmd_beat_count = 3'h0;
  end
  if (reset) begin
    ifu_bus_arready_unq_ff = 1'h0;
  end
  if (reset) begin
    ifu_bus_arvalid_ff = 1'h0;
  end
  if (reset) begin
    ifc_dma_access_ok_prev = 1'h0;
  end
  if (reset) begin
    iccm_ecc_corr_data_ff = 39'h0;
  end
  if (reset) begin
    dma_mem_addr_ff = 2'h0;
  end
  if (reset) begin
    dma_mem_tag_ff = 3'h0;
  end
  if (reset) begin
    iccm_dma_rtag_temp = 3'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_temp = 1'h0;
  end
  if (reset) begin
    iccm_dma_ecc_error = 1'h0;
  end
  if (reset) begin
    iccm_dma_rdata_temp = 64'h0;
  end
  if (reset) begin
    iccm_ecc_corr_index_ff = 14'h0;
  end
  if (reset) begin
    iccm_rd_ecc_single_err_ff = 1'h0;
  end
  if (reset) begin
    iccm_rw_addr_f = 14'h0;
  end
  if (reset) begin
    ifu_status_wr_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_wr_en_ff = 1'h0;
  end
  if (reset) begin
    way_status_new_ff = 1'h0;
  end
  if (reset) begin
    ifu_tag_wren_ff = 2'h0;
  end
  if (reset) begin
    ic_valid_ff = 1'h0;
  end
  if (reset) begin
    _T_10552 = 1'h0;
  end
  if (reset) begin
    _T_10556 = 1'h0;
  end
  if (reset) begin
    _T_10561 = 1'h0;
  end
  if (reset) begin
    _T_10568 = 1'h0;
  end
  if (reset) begin
    _T_10572 = 1'h0;
  end
  if (reset) begin
    _T_10598 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else if (_T_1) begin
      flush_final_f <= io_exu_flush_final;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else if (_T_337) begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_27) begin
        if (_T_29) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_34) begin
        if (_T_39) begin
          miss_state <= 3'h0;
        end else if (_T_43) begin
          miss_state <= 3'h3;
        end else if (_T_50) begin
          miss_state <= 3'h4;
        end else if (_T_54) begin
          miss_state <= 3'h0;
        end else if (_T_64) begin
          miss_state <= 3'h6;
        end else if (_T_74) begin
          miss_state <= 3'h6;
        end else if (_T_82) begin
          miss_state <= 3'h0;
        end else if (_T_87) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_105) begin
        miss_state <= 3'h0;
      end else if (_T_109) begin
        if (_T_116) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_124) begin
        if (_T_129) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_135) begin
        if (_T_140) begin
          miss_state <= 3'h5;
        end else if (_T_146) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_154) begin
        if (io_dec_mem_ctrl_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_35) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_163) begin
        if (io_dec_mem_ctrl_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_35) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else if (_T_2613) begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else if (fetch_bf_f_c1_clken) begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else if (fetch_bf_f_c1_clken) begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else if (_T_3169) begin
      iccm_dma_rvalid_in <= _T_2764;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else if (_T_2757) begin
      dma_iccm_req_f <= io_dma_mem_ctl_dma_iccm_req;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2521) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2523) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2533) begin
        perr_state <= 3'h0;
      end else if (_T_2536) begin
        if (_T_2539) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2543) begin
        if (io_dec_mem_ctrl_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2547) begin
        err_stop_state <= 2'h1;
      end else if (_T_2552) begin
        if (_T_2554) begin
          err_stop_state <= 2'h0;
        end else if (_T_2575) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2579) begin
        if (_T_2554) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2596) begin
        if (_T_2600) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_mem_ctrl_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else if (_T_4081) begin
      reset_all_tags <= io_dec_mem_ctrl_dec_tlu_fence_i_wb;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else if (fetch_bf_f_c1_clken) begin
      ifc_region_acc_fault_final_f <= ifc_region_acc_fault_final_bf;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_r_valid;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else if (_T_2609) begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (fetch_bf_f_c1_clken) begin
      if (scnd_miss_req) begin
        uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
      end else if (!(sel_hold_imb)) begin
        uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else if (_T_2668) begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= {_T_1390,ic_miss_buff_data_valid_in_0};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      imb_ff <= 31'h0;
    end else if (fetch_bf_f_c1_clken) begin
      if (scnd_miss_req) begin
        imb_ff <= imb_scnd_ff;
      end else if (!(sel_hold_imb)) begin
        imb_ff <= io_ifc_fetch_addr_bf;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else if (_T_2677) begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else if (_T_375) begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (fetch_bf_f_c1_clken) begin
      if (!(_T_22)) begin
        way_status_mb_scnd_ff <= way_status;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_5290) begin
      if (_T_4089) begin
        ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
      end else begin
        ifu_ic_rw_int_addr_ff <= io_ic_rw_addr[11:5];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_4123) begin
      way_status_out_0 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_4128) begin
      way_status_out_1 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_4133) begin
      way_status_out_2 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_4138) begin
      way_status_out_3 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_4143) begin
      way_status_out_4 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_4148) begin
      way_status_out_5 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_4153) begin
      way_status_out_6 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_4158) begin
      way_status_out_7 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_4163) begin
      way_status_out_8 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_4168) begin
      way_status_out_9 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_4173) begin
      way_status_out_10 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_4178) begin
      way_status_out_11 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_4183) begin
      way_status_out_12 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_4188) begin
      way_status_out_13 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_4193) begin
      way_status_out_14 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_4198) begin
      way_status_out_15 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_4203) begin
      way_status_out_16 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_4208) begin
      way_status_out_17 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_4213) begin
      way_status_out_18 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_4218) begin
      way_status_out_19 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_4223) begin
      way_status_out_20 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_4228) begin
      way_status_out_21 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_4233) begin
      way_status_out_22 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_4238) begin
      way_status_out_23 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_4243) begin
      way_status_out_24 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_4248) begin
      way_status_out_25 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_4253) begin
      way_status_out_26 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_4258) begin
      way_status_out_27 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_4263) begin
      way_status_out_28 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_4268) begin
      way_status_out_29 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_4273) begin
      way_status_out_30 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_4278) begin
      way_status_out_31 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_4283) begin
      way_status_out_32 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_4288) begin
      way_status_out_33 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_4293) begin
      way_status_out_34 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_4298) begin
      way_status_out_35 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_4303) begin
      way_status_out_36 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_4308) begin
      way_status_out_37 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_4313) begin
      way_status_out_38 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_4318) begin
      way_status_out_39 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_4323) begin
      way_status_out_40 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_4328) begin
      way_status_out_41 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_4333) begin
      way_status_out_42 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_4338) begin
      way_status_out_43 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_4343) begin
      way_status_out_44 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_4348) begin
      way_status_out_45 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_4353) begin
      way_status_out_46 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_4358) begin
      way_status_out_47 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_4363) begin
      way_status_out_48 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_4368) begin
      way_status_out_49 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_4373) begin
      way_status_out_50 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_4378) begin
      way_status_out_51 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_4383) begin
      way_status_out_52 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_4388) begin
      way_status_out_53 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_4393) begin
      way_status_out_54 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_4398) begin
      way_status_out_55 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_4403) begin
      way_status_out_56 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_4408) begin
      way_status_out_57 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_4413) begin
      way_status_out_58 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_4418) begin
      way_status_out_59 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_4423) begin
      way_status_out_60 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_4428) begin
      way_status_out_61 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_4433) begin
      way_status_out_62 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_4438) begin
      way_status_out_63 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_4443) begin
      way_status_out_64 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_4448) begin
      way_status_out_65 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_4453) begin
      way_status_out_66 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_4458) begin
      way_status_out_67 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_4463) begin
      way_status_out_68 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_4468) begin
      way_status_out_69 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_4473) begin
      way_status_out_70 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_4478) begin
      way_status_out_71 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_4483) begin
      way_status_out_72 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_4488) begin
      way_status_out_73 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_4493) begin
      way_status_out_74 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_4498) begin
      way_status_out_75 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_4503) begin
      way_status_out_76 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_4508) begin
      way_status_out_77 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_4513) begin
      way_status_out_78 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_4518) begin
      way_status_out_79 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_4523) begin
      way_status_out_80 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_4528) begin
      way_status_out_81 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_4533) begin
      way_status_out_82 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_4538) begin
      way_status_out_83 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_4543) begin
      way_status_out_84 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_4548) begin
      way_status_out_85 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_4553) begin
      way_status_out_86 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_4558) begin
      way_status_out_87 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_4563) begin
      way_status_out_88 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_4568) begin
      way_status_out_89 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_4573) begin
      way_status_out_90 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_4578) begin
      way_status_out_91 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_4583) begin
      way_status_out_92 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_4588) begin
      way_status_out_93 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_4593) begin
      way_status_out_94 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_4598) begin
      way_status_out_95 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_4603) begin
      way_status_out_96 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_4608) begin
      way_status_out_97 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_4613) begin
      way_status_out_98 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_4618) begin
      way_status_out_99 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_4623) begin
      way_status_out_100 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_4628) begin
      way_status_out_101 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_4633) begin
      way_status_out_102 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_4638) begin
      way_status_out_103 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_4643) begin
      way_status_out_104 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_4648) begin
      way_status_out_105 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_4653) begin
      way_status_out_106 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_4658) begin
      way_status_out_107 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_4663) begin
      way_status_out_108 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_4668) begin
      way_status_out_109 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_4673) begin
      way_status_out_110 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_4678) begin
      way_status_out_111 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_4683) begin
      way_status_out_112 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_4688) begin
      way_status_out_113 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_4693) begin
      way_status_out_114 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_4698) begin
      way_status_out_115 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_4703) begin
      way_status_out_116 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_4708) begin
      way_status_out_117 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_4713) begin
      way_status_out_118 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_4718) begin
      way_status_out_119 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_4723) begin
      way_status_out_120 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_4728) begin
      way_status_out_121 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_4733) begin
      way_status_out_122 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_4738) begin
      way_status_out_123 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_4743) begin
      way_status_out_124 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_4748) begin
      way_status_out_125 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_4753) begin
      way_status_out_126 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_4758) begin
      way_status_out_127 <= way_status_new_ff;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      tagv_mb_scnd_ff <= 2'h0;
    end else if (fetch_bf_f_c1_clken) begin
      if (!(_T_22)) begin
        tagv_mb_scnd_ff <= _T_203;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (fetch_bf_f_c1_clken) begin
      if (!(sel_hold_imb_scnd)) begin
        uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (fetch_bf_f_c1_clken) begin
      if (!(sel_hold_imb_scnd)) begin
        imb_scnd_ff <= io_ifc_fetch_addr_bf;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_r_bits_id;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_r_bits_resp;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else if (_T_1272) begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (fetch_bf_f_c1_clken) begin
      if (_T_284) begin
        way_status_mb_ff <= way_status_mb_scnd_ff;
      end else if (_T_286) begin
        way_status_mb_ff <= replace_way_mb_any_0;
      end else if (!(miss_pending)) begin
        way_status_mb_ff <= way_status;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (fetch_bf_f_c1_clken) begin
      if (scnd_miss_req) begin
        tagv_mb_ff <= _T_296;
      end else if (!(miss_pending)) begin
        tagv_mb_ff <= _T_303;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      reset_ic_ff <= 1'h0;
    end else if (_T_310) begin
      reset_ic_ff <= reset_ic_in;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else if (_T_313) begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_326) begin
      if (_T_237) begin
        miss_addr <= imb_ff[30:5];
      end else if (scnd_miss_req_q) begin
        miss_addr <= imb_scnd_ff[30:5];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else if (fetch_bf_f_c1_clken) begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_326) begin
      if (_T_237) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2683;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else if (_T_2728) begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (_T_377) begin
      ifu_bus_rdata_ff <= io_ifu_axi_r_bits_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else if (_T_1554) begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= {_T_1430,ic_miss_buff_data_error_in_0};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5947) begin
      ic_tag_valid_out_1_0 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5964) begin
      ic_tag_valid_out_1_1 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5981) begin
      ic_tag_valid_out_1_2 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5998) begin
      ic_tag_valid_out_1_3 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_6015) begin
      ic_tag_valid_out_1_4 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_6032) begin
      ic_tag_valid_out_1_5 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_6049) begin
      ic_tag_valid_out_1_6 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_6066) begin
      ic_tag_valid_out_1_7 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_6083) begin
      ic_tag_valid_out_1_8 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_6100) begin
      ic_tag_valid_out_1_9 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_6117) begin
      ic_tag_valid_out_1_10 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_6134) begin
      ic_tag_valid_out_1_11 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_6151) begin
      ic_tag_valid_out_1_12 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_6168) begin
      ic_tag_valid_out_1_13 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_6185) begin
      ic_tag_valid_out_1_14 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_6202) begin
      ic_tag_valid_out_1_15 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_6219) begin
      ic_tag_valid_out_1_16 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_6236) begin
      ic_tag_valid_out_1_17 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_6253) begin
      ic_tag_valid_out_1_18 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_6270) begin
      ic_tag_valid_out_1_19 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_6287) begin
      ic_tag_valid_out_1_20 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_6304) begin
      ic_tag_valid_out_1_21 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_6321) begin
      ic_tag_valid_out_1_22 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_6338) begin
      ic_tag_valid_out_1_23 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6355) begin
      ic_tag_valid_out_1_24 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6372) begin
      ic_tag_valid_out_1_25 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6389) begin
      ic_tag_valid_out_1_26 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6406) begin
      ic_tag_valid_out_1_27 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6423) begin
      ic_tag_valid_out_1_28 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6440) begin
      ic_tag_valid_out_1_29 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6457) begin
      ic_tag_valid_out_1_30 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6474) begin
      ic_tag_valid_out_1_31 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_7035) begin
      ic_tag_valid_out_1_32 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_7052) begin
      ic_tag_valid_out_1_33 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_7069) begin
      ic_tag_valid_out_1_34 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_7086) begin
      ic_tag_valid_out_1_35 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_7103) begin
      ic_tag_valid_out_1_36 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_7120) begin
      ic_tag_valid_out_1_37 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_7137) begin
      ic_tag_valid_out_1_38 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_7154) begin
      ic_tag_valid_out_1_39 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_7171) begin
      ic_tag_valid_out_1_40 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_7188) begin
      ic_tag_valid_out_1_41 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_7205) begin
      ic_tag_valid_out_1_42 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_7222) begin
      ic_tag_valid_out_1_43 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_7239) begin
      ic_tag_valid_out_1_44 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_7256) begin
      ic_tag_valid_out_1_45 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_7273) begin
      ic_tag_valid_out_1_46 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_7290) begin
      ic_tag_valid_out_1_47 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_7307) begin
      ic_tag_valid_out_1_48 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_7324) begin
      ic_tag_valid_out_1_49 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_7341) begin
      ic_tag_valid_out_1_50 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_7358) begin
      ic_tag_valid_out_1_51 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_7375) begin
      ic_tag_valid_out_1_52 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_7392) begin
      ic_tag_valid_out_1_53 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_7409) begin
      ic_tag_valid_out_1_54 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_7426) begin
      ic_tag_valid_out_1_55 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_7443) begin
      ic_tag_valid_out_1_56 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_7460) begin
      ic_tag_valid_out_1_57 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_7477) begin
      ic_tag_valid_out_1_58 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7494) begin
      ic_tag_valid_out_1_59 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7511) begin
      ic_tag_valid_out_1_60 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7528) begin
      ic_tag_valid_out_1_61 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7545) begin
      ic_tag_valid_out_1_62 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7562) begin
      ic_tag_valid_out_1_63 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_8123) begin
      ic_tag_valid_out_1_64 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_8140) begin
      ic_tag_valid_out_1_65 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_8157) begin
      ic_tag_valid_out_1_66 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_8174) begin
      ic_tag_valid_out_1_67 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_8191) begin
      ic_tag_valid_out_1_68 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_8208) begin
      ic_tag_valid_out_1_69 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_8225) begin
      ic_tag_valid_out_1_70 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_8242) begin
      ic_tag_valid_out_1_71 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_8259) begin
      ic_tag_valid_out_1_72 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_8276) begin
      ic_tag_valid_out_1_73 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_8293) begin
      ic_tag_valid_out_1_74 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_8310) begin
      ic_tag_valid_out_1_75 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_8327) begin
      ic_tag_valid_out_1_76 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_8344) begin
      ic_tag_valid_out_1_77 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_8361) begin
      ic_tag_valid_out_1_78 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_8378) begin
      ic_tag_valid_out_1_79 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_8395) begin
      ic_tag_valid_out_1_80 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_8412) begin
      ic_tag_valid_out_1_81 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_8429) begin
      ic_tag_valid_out_1_82 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_8446) begin
      ic_tag_valid_out_1_83 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_8463) begin
      ic_tag_valid_out_1_84 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_8480) begin
      ic_tag_valid_out_1_85 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_8497) begin
      ic_tag_valid_out_1_86 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_8514) begin
      ic_tag_valid_out_1_87 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8531) begin
      ic_tag_valid_out_1_88 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8548) begin
      ic_tag_valid_out_1_89 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8565) begin
      ic_tag_valid_out_1_90 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8582) begin
      ic_tag_valid_out_1_91 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8599) begin
      ic_tag_valid_out_1_92 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8616) begin
      ic_tag_valid_out_1_93 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8633) begin
      ic_tag_valid_out_1_94 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8650) begin
      ic_tag_valid_out_1_95 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_9211) begin
      ic_tag_valid_out_1_96 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_9228) begin
      ic_tag_valid_out_1_97 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_9245) begin
      ic_tag_valid_out_1_98 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_9262) begin
      ic_tag_valid_out_1_99 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_9279) begin
      ic_tag_valid_out_1_100 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_9296) begin
      ic_tag_valid_out_1_101 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_9313) begin
      ic_tag_valid_out_1_102 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_9330) begin
      ic_tag_valid_out_1_103 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_9347) begin
      ic_tag_valid_out_1_104 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_9364) begin
      ic_tag_valid_out_1_105 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_9381) begin
      ic_tag_valid_out_1_106 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_9398) begin
      ic_tag_valid_out_1_107 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_9415) begin
      ic_tag_valid_out_1_108 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_9432) begin
      ic_tag_valid_out_1_109 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_9449) begin
      ic_tag_valid_out_1_110 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_9466) begin
      ic_tag_valid_out_1_111 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_9483) begin
      ic_tag_valid_out_1_112 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_9500) begin
      ic_tag_valid_out_1_113 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_9517) begin
      ic_tag_valid_out_1_114 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9534) begin
      ic_tag_valid_out_1_115 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9551) begin
      ic_tag_valid_out_1_116 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9568) begin
      ic_tag_valid_out_1_117 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9585) begin
      ic_tag_valid_out_1_118 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9602) begin
      ic_tag_valid_out_1_119 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_9619) begin
      ic_tag_valid_out_1_120 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_9636) begin
      ic_tag_valid_out_1_121 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_9653) begin
      ic_tag_valid_out_1_122 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_9670) begin
      ic_tag_valid_out_1_123 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_9687) begin
      ic_tag_valid_out_1_124 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_9704) begin
      ic_tag_valid_out_1_125 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_9721) begin
      ic_tag_valid_out_1_126 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_9738) begin
      ic_tag_valid_out_1_127 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5403) begin
      ic_tag_valid_out_0_0 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5420) begin
      ic_tag_valid_out_0_1 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5437) begin
      ic_tag_valid_out_0_2 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5454) begin
      ic_tag_valid_out_0_3 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5471) begin
      ic_tag_valid_out_0_4 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5488) begin
      ic_tag_valid_out_0_5 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5505) begin
      ic_tag_valid_out_0_6 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5522) begin
      ic_tag_valid_out_0_7 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5539) begin
      ic_tag_valid_out_0_8 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5556) begin
      ic_tag_valid_out_0_9 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5573) begin
      ic_tag_valid_out_0_10 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5590) begin
      ic_tag_valid_out_0_11 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5607) begin
      ic_tag_valid_out_0_12 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5624) begin
      ic_tag_valid_out_0_13 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5641) begin
      ic_tag_valid_out_0_14 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5658) begin
      ic_tag_valid_out_0_15 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5675) begin
      ic_tag_valid_out_0_16 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5692) begin
      ic_tag_valid_out_0_17 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5709) begin
      ic_tag_valid_out_0_18 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5726) begin
      ic_tag_valid_out_0_19 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5743) begin
      ic_tag_valid_out_0_20 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5760) begin
      ic_tag_valid_out_0_21 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5777) begin
      ic_tag_valid_out_0_22 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5794) begin
      ic_tag_valid_out_0_23 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5811) begin
      ic_tag_valid_out_0_24 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5828) begin
      ic_tag_valid_out_0_25 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5845) begin
      ic_tag_valid_out_0_26 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5862) begin
      ic_tag_valid_out_0_27 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5879) begin
      ic_tag_valid_out_0_28 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5896) begin
      ic_tag_valid_out_0_29 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5913) begin
      ic_tag_valid_out_0_30 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5930) begin
      ic_tag_valid_out_0_31 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6491) begin
      ic_tag_valid_out_0_32 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6508) begin
      ic_tag_valid_out_0_33 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6525) begin
      ic_tag_valid_out_0_34 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6542) begin
      ic_tag_valid_out_0_35 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6559) begin
      ic_tag_valid_out_0_36 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6576) begin
      ic_tag_valid_out_0_37 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6593) begin
      ic_tag_valid_out_0_38 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6610) begin
      ic_tag_valid_out_0_39 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6627) begin
      ic_tag_valid_out_0_40 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6644) begin
      ic_tag_valid_out_0_41 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6661) begin
      ic_tag_valid_out_0_42 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6678) begin
      ic_tag_valid_out_0_43 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6695) begin
      ic_tag_valid_out_0_44 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6712) begin
      ic_tag_valid_out_0_45 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6729) begin
      ic_tag_valid_out_0_46 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6746) begin
      ic_tag_valid_out_0_47 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6763) begin
      ic_tag_valid_out_0_48 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6780) begin
      ic_tag_valid_out_0_49 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6797) begin
      ic_tag_valid_out_0_50 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6814) begin
      ic_tag_valid_out_0_51 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6831) begin
      ic_tag_valid_out_0_52 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6848) begin
      ic_tag_valid_out_0_53 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6865) begin
      ic_tag_valid_out_0_54 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6882) begin
      ic_tag_valid_out_0_55 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6899) begin
      ic_tag_valid_out_0_56 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6916) begin
      ic_tag_valid_out_0_57 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6933) begin
      ic_tag_valid_out_0_58 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6950) begin
      ic_tag_valid_out_0_59 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6967) begin
      ic_tag_valid_out_0_60 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6984) begin
      ic_tag_valid_out_0_61 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_7001) begin
      ic_tag_valid_out_0_62 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_7018) begin
      ic_tag_valid_out_0_63 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7579) begin
      ic_tag_valid_out_0_64 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7596) begin
      ic_tag_valid_out_0_65 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7613) begin
      ic_tag_valid_out_0_66 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7630) begin
      ic_tag_valid_out_0_67 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7647) begin
      ic_tag_valid_out_0_68 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7664) begin
      ic_tag_valid_out_0_69 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7681) begin
      ic_tag_valid_out_0_70 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7698) begin
      ic_tag_valid_out_0_71 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7715) begin
      ic_tag_valid_out_0_72 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7732) begin
      ic_tag_valid_out_0_73 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7749) begin
      ic_tag_valid_out_0_74 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7766) begin
      ic_tag_valid_out_0_75 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7783) begin
      ic_tag_valid_out_0_76 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7800) begin
      ic_tag_valid_out_0_77 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7817) begin
      ic_tag_valid_out_0_78 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7834) begin
      ic_tag_valid_out_0_79 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7851) begin
      ic_tag_valid_out_0_80 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7868) begin
      ic_tag_valid_out_0_81 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7885) begin
      ic_tag_valid_out_0_82 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7902) begin
      ic_tag_valid_out_0_83 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7919) begin
      ic_tag_valid_out_0_84 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7936) begin
      ic_tag_valid_out_0_85 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7953) begin
      ic_tag_valid_out_0_86 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7970) begin
      ic_tag_valid_out_0_87 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7987) begin
      ic_tag_valid_out_0_88 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_8004) begin
      ic_tag_valid_out_0_89 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_8021) begin
      ic_tag_valid_out_0_90 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_8038) begin
      ic_tag_valid_out_0_91 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_8055) begin
      ic_tag_valid_out_0_92 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_8072) begin
      ic_tag_valid_out_0_93 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_8089) begin
      ic_tag_valid_out_0_94 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_8106) begin
      ic_tag_valid_out_0_95 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8667) begin
      ic_tag_valid_out_0_96 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8684) begin
      ic_tag_valid_out_0_97 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8701) begin
      ic_tag_valid_out_0_98 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8718) begin
      ic_tag_valid_out_0_99 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8735) begin
      ic_tag_valid_out_0_100 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8752) begin
      ic_tag_valid_out_0_101 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8769) begin
      ic_tag_valid_out_0_102 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8786) begin
      ic_tag_valid_out_0_103 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8803) begin
      ic_tag_valid_out_0_104 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8820) begin
      ic_tag_valid_out_0_105 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8837) begin
      ic_tag_valid_out_0_106 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8854) begin
      ic_tag_valid_out_0_107 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8871) begin
      ic_tag_valid_out_0_108 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8888) begin
      ic_tag_valid_out_0_109 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8905) begin
      ic_tag_valid_out_0_110 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8922) begin
      ic_tag_valid_out_0_111 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8939) begin
      ic_tag_valid_out_0_112 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8956) begin
      ic_tag_valid_out_0_113 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8973) begin
      ic_tag_valid_out_0_114 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8990) begin
      ic_tag_valid_out_0_115 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_9007) begin
      ic_tag_valid_out_0_116 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_9024) begin
      ic_tag_valid_out_0_117 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_9041) begin
      ic_tag_valid_out_0_118 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_9058) begin
      ic_tag_valid_out_0_119 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_9075) begin
      ic_tag_valid_out_0_120 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_9092) begin
      ic_tag_valid_out_0_121 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_9109) begin
      ic_tag_valid_out_0_122 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_9126) begin
      ic_tag_valid_out_0_123 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_9143) begin
      ic_tag_valid_out_0_124 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_9160) begin
      ic_tag_valid_out_0_125 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_9177) begin
      ic_tag_valid_out_0_126 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_9194) begin
      ic_tag_valid_out_0_127 <= _T_5392;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else if (_T_10593) begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1237 <= 71'h0;
    end else if (ic_debug_rd_en_ff) begin
      if (ic_debug_ict_array_sel_ff) begin
        _T_1237 <= _T_1236;
      end else begin
        _T_1237 <= io_ic_debug_rd_data;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_memory_f <= 1'h0;
    end else if (_T_10661) begin
      ifc_region_acc_fault_memory_f <= ifc_region_acc_fault_memory_bf;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else if (_T_2517) begin
      dma_sb_err_state_ff <= _T_10;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      bus_cmd_req_hold <= 1'h0;
    end else if (_T_2635) begin
      bus_cmd_req_hold <= bus_cmd_req_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2627) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2711) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_ar_ready;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_ar_valid;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else if (_T_2744) begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_4021;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else if (_T_3166) begin
      dma_mem_addr_ff <= io_dma_mem_ctl_dma_mem_addr[3:2];
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else if (_T_3158) begin
      dma_mem_tag_ff <= io_dma_mem_ctl_dma_mem_tag;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rtag_temp <= 3'h0;
    end else if (_T_3161) begin
      iccm_dma_rtag_temp <= dma_mem_tag_ff;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_temp <= 1'h0;
    end else if (_T_3172) begin
      iccm_dma_rvalid_temp <= iccm_dma_rvalid_in;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      iccm_dma_ecc_error <= 1'h0;
    end else if (_T_3176) begin
      iccm_dma_ecc_error <= _T_3154;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      iccm_dma_rdata_temp <= 64'h0;
    end else if (iccm_dma_rvalid_in) begin
      if (_T_3154) begin
        iccm_dma_rdata_temp <= _T_3155;
      end else begin
        iccm_dma_rdata_temp <= _T_3156;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_4015;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else if (_T_4003) begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else if (_T_4019) begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_4093) begin
      if (_T_4089) begin
        ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
      end else begin
        ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else if (_T_4097) begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_4102) begin
      if (_T_4095) begin
        way_status_new_ff <= io_ic_debug_wr_data[4];
      end else if (_T_10527) begin
        way_status_new_ff <= replace_way_mb_any_0;
      end else begin
        way_status_new_ff <= way_status_hit_new;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else if (_T_5293) begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_5298) begin
      if (_T_4095) begin
        ic_valid_ff <= io_ic_debug_wr_data[0];
      end else begin
        ic_valid_ff <= ic_valid;
      end
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      _T_10552 <= 1'h0;
    end else if (_T_10551) begin
      _T_10552 <= ic_act_miss_f;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      _T_10556 <= 1'h0;
    end else if (_T_10555) begin
      _T_10556 <= ic_act_hit_f;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      _T_10561 <= 1'h0;
    end else if (_T_10560) begin
      _T_10561 <= _T_2500;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      _T_10568 <= 1'h0;
    end else if (_T_10567) begin
      _T_10568 <= _T_10564;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      _T_10572 <= 1'h0;
    end else if (_T_10571) begin
      _T_10572 <= bus_cmd_sent;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      _T_10598 <= 1'h0;
    end else if (_T_10597) begin
      _T_10598 <= ic_debug_rd_en_ff;
    end
  end
endmodule
module ifu_bp_ctl(
  input         clock,
  input         reset,
  input         io_ic_hit_f,
  input         io_exu_flush_final,
  input  [30:0] io_ifc_fetch_addr_f,
  input         io_ifc_fetch_req_f,
  input         io_dec_bp_dec_tlu_br0_r_pkt_valid,
  input  [1:0]  io_dec_bp_dec_tlu_br0_r_pkt_bits_hist,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_way,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_middle,
  input         io_dec_bp_dec_tlu_flush_leak_one_wb,
  input         io_dec_bp_dec_tlu_bpred_disable,
  input         io_dec_tlu_flush_lower_wb,
  input  [7:0]  io_exu_bp_exu_i0_br_index_r,
  input  [7:0]  io_exu_bp_exu_i0_br_fghr_r,
  input         io_exu_bp_exu_mp_pkt_valid,
  input         io_exu_bp_exu_mp_pkt_bits_misp,
  input         io_exu_bp_exu_mp_pkt_bits_ataken,
  input         io_exu_bp_exu_mp_pkt_bits_boffset,
  input         io_exu_bp_exu_mp_pkt_bits_pc4,
  input  [1:0]  io_exu_bp_exu_mp_pkt_bits_hist,
  input  [11:0] io_exu_bp_exu_mp_pkt_bits_toffset,
  input         io_exu_bp_exu_mp_pkt_bits_pcall,
  input         io_exu_bp_exu_mp_pkt_bits_pja,
  input         io_exu_bp_exu_mp_pkt_bits_way,
  input         io_exu_bp_exu_mp_pkt_bits_pret,
  input  [7:0]  io_exu_bp_exu_mp_eghr,
  input  [7:0]  io_exu_bp_exu_mp_fghr,
  input  [7:0]  io_exu_bp_exu_mp_index,
  input  [4:0]  io_exu_bp_exu_mp_btag,
  output        io_ifu_bp_hit_taken_f,
  output [30:0] io_ifu_bp_btb_target_f,
  output        io_ifu_bp_inst_mask_f,
  output [7:0]  io_ifu_bp_fghr_f,
  output [1:0]  io_ifu_bp_way_f,
  output [1:0]  io_ifu_bp_ret_f,
  output [1:0]  io_ifu_bp_hist1_f,
  output [1:0]  io_ifu_bp_hist0_f,
  output [1:0]  io_ifu_bp_pc4_f,
  output [1:0]  io_ifu_bp_valid_f,
  output [11:0] io_ifu_bp_poffset_f
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [255:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_13_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_14_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_15_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_16_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_17_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_18_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_19_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_20_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_20_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_21_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_21_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_22_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_22_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_23_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_23_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_24_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_24_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_25_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_25_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_26_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_26_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_27_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_27_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_28_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_28_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_29_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_29_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_30_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_30_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_31_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_31_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_32_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_32_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_33_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_33_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_34_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_34_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_35_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_35_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_36_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_36_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_37_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_37_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_38_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_38_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_39_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_39_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_40_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_40_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_41_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_41_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_42_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_42_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_43_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_43_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_44_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_44_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_45_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_45_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_46_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_46_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_47_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_47_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_48_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_48_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_49_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_49_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_50_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_50_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_51_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_51_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_52_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_52_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_53_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_53_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_54_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_54_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_55_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_55_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_56_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_56_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_57_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_57_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_58_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_58_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_59_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_59_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_60_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_60_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_61_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_61_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_62_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_62_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_63_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_63_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_64_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_64_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_65_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_65_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_66_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_66_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_67_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_67_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_68_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_68_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_69_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_69_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_70_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_70_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_71_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_71_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_72_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_72_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_73_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_73_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_74_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_74_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_75_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_75_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_76_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_76_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_77_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_77_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_78_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_78_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_79_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_79_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_80_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_80_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_81_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_81_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_82_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_82_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_83_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_83_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_84_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_84_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_85_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_85_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_86_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_86_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_87_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_87_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_88_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_88_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_89_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_89_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_90_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_90_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_91_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_91_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_92_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_92_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_93_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_93_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_94_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_94_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_95_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_95_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_96_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_96_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_97_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_97_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_98_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_98_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_99_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_99_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_100_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_100_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_101_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_101_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_102_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_102_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_103_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_103_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_104_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_104_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_105_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_105_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_106_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_106_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_107_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_107_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_108_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_108_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_109_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_109_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_110_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_110_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_111_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_111_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_112_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_112_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_113_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_113_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_114_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_114_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_115_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_115_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_116_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_116_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_117_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_117_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_118_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_118_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_119_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_119_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_120_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_120_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_121_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_121_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_122_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_122_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_123_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_123_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_124_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_124_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_125_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_125_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_126_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_126_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_127_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_127_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_128_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_128_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_129_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_129_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_130_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_130_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_131_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_131_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_132_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_132_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_133_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_133_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_134_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_134_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_135_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_135_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_136_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_136_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_137_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_137_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_138_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_138_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_139_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_139_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_140_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_140_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_141_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_141_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_142_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_142_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_143_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_143_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_144_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_144_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_145_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_145_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_146_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_146_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_147_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_147_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_148_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_148_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_149_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_149_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_150_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_150_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_151_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_151_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_152_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_152_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_153_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_153_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_154_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_154_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_155_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_155_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_156_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_156_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_157_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_157_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_158_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_158_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_159_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_159_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_160_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_160_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_161_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_161_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_162_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_162_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_163_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_163_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_164_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_164_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_165_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_165_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_166_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_166_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_167_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_167_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_168_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_168_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_169_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_169_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_170_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_170_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_171_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_171_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_172_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_172_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_173_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_173_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_174_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_174_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_175_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_175_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_176_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_176_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_177_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_177_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_178_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_178_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_179_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_179_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_180_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_180_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_181_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_181_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_182_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_182_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_183_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_183_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_184_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_184_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_185_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_185_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_186_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_186_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_187_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_187_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_188_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_188_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_189_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_189_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_190_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_190_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_191_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_191_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_192_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_192_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_193_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_193_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_194_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_194_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_195_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_195_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_196_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_196_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_197_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_197_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_198_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_198_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_199_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_199_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_200_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_200_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_201_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_201_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_202_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_202_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_203_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_203_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_204_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_204_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_205_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_205_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_206_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_206_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_207_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_207_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_208_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_208_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_209_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_209_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_210_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_210_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_211_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_211_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_212_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_212_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_213_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_213_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_214_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_214_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_215_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_215_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_216_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_216_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_217_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_217_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_218_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_218_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_219_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_219_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_220_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_220_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_221_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_221_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_222_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_222_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_223_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_223_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_224_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_224_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_225_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_225_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_226_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_226_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_227_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_227_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_228_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_228_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_229_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_229_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_230_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_230_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_231_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_231_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_232_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_232_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_233_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_233_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_234_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_234_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_235_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_235_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_236_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_236_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_237_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_237_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_238_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_238_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_239_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_239_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_240_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_240_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_241_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_241_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_242_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_242_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_243_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_243_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_244_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_244_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_245_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_245_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_246_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_246_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_247_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_247_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_248_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_248_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_249_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_249_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_250_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_250_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_251_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_251_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_252_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_252_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_253_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_253_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_254_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_254_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_255_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_255_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_256_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_256_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_257_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_257_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_258_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_258_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_259_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_259_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_260_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_260_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_261_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_261_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_262_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_262_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_263_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_263_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_264_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_264_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_265_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_265_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_266_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_266_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_267_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_267_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_268_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_268_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_269_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_269_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_270_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_270_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_271_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_271_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_272_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_272_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_273_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_273_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_274_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_274_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_275_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_275_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_276_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_276_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_277_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_277_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_278_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_278_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_279_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_279_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_280_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_280_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_281_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_281_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_282_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_282_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_283_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_283_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_284_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_284_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_285_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_285_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_286_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_286_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_287_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_287_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_288_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_288_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_289_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_289_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_290_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_290_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_291_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_291_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_292_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_292_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_293_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_293_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_294_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_294_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_295_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_295_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_296_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_296_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_297_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_297_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_298_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_298_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_299_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_299_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_300_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_300_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_301_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_301_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_302_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_302_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_303_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_303_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_304_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_304_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_305_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_305_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_306_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_306_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_307_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_307_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_308_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_308_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_309_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_309_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_310_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_310_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_311_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_311_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_312_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_312_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_313_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_313_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_314_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_314_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_315_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_315_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_316_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_316_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_317_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_317_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_318_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_318_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_319_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_319_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_320_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_320_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_321_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_321_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_322_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_322_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_323_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_323_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_324_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_324_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_325_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_325_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_326_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_326_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_327_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_327_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_328_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_328_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_329_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_329_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_330_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_330_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_331_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_331_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_332_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_332_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_333_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_333_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_334_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_334_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_335_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_335_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_336_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_336_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_337_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_337_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_338_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_338_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_339_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_339_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_340_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_340_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_341_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_341_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_342_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_342_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_343_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_343_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_344_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_344_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_345_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_345_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_346_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_346_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_347_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_347_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_348_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_348_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_349_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_349_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_350_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_350_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_351_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_351_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_352_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_352_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_353_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_353_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_354_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_354_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_355_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_355_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_356_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_356_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_357_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_357_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_358_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_358_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_359_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_359_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_360_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_360_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_361_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_361_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_362_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_362_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_363_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_363_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_364_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_364_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_365_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_365_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_366_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_366_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_367_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_367_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_368_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_368_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_369_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_369_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_370_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_370_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_371_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_371_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_372_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_372_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_373_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_373_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_374_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_374_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_375_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_375_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_376_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_376_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_377_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_377_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_378_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_378_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_379_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_379_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_380_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_380_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_381_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_381_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_382_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_382_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_383_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_383_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_384_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_384_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_385_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_385_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_386_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_386_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_387_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_387_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_388_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_388_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_389_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_389_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_390_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_390_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_391_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_391_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_392_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_392_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_393_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_393_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_394_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_394_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_395_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_395_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_396_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_396_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_397_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_397_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_398_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_398_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_399_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_399_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_400_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_400_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_401_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_401_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_402_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_402_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_403_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_403_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_404_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_404_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_405_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_405_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_406_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_406_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_407_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_407_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_408_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_408_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_409_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_409_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_410_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_410_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_411_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_411_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_412_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_412_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_413_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_413_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_414_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_414_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_415_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_415_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_416_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_416_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_417_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_417_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_418_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_418_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_419_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_419_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_420_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_420_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_421_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_421_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_422_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_422_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_423_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_423_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_424_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_424_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_425_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_425_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_426_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_426_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_427_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_427_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_428_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_428_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_429_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_429_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_430_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_430_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_431_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_431_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_432_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_432_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_433_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_433_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_434_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_434_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_435_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_435_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_436_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_436_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_437_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_437_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_438_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_438_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_439_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_439_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_440_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_440_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_441_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_441_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_442_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_442_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_443_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_443_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_444_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_444_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_445_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_445_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_446_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_446_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_447_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_447_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_448_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_448_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_449_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_449_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_450_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_450_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_451_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_451_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_452_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_452_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_453_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_453_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_454_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_454_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_455_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_455_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_456_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_456_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_457_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_457_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_458_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_458_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_459_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_459_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_460_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_460_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_461_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_461_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_462_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_462_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_463_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_463_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_464_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_464_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_465_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_465_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_466_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_466_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_467_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_467_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_468_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_468_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_469_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_469_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_470_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_470_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_471_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_471_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_472_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_472_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_473_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_473_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_474_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_474_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_475_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_475_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_476_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_476_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_477_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_477_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_478_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_478_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_479_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_479_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_480_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_480_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_481_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_481_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_482_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_482_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_483_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_483_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_484_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_484_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_485_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_485_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_486_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_486_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_487_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_487_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_488_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_488_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_489_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_489_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_490_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_490_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_491_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_491_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_492_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_492_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_493_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_493_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_494_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_494_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_495_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_495_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_496_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_496_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_497_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_497_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_498_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_498_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_499_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_499_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_500_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_500_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_501_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_501_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_502_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_502_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_503_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_503_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_504_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_504_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_505_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_505_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_506_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_506_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_507_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_507_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_508_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_508_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_509_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_509_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_510_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_510_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_511_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_511_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_512_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_512_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_513_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_513_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_514_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_514_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_515_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_515_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_516_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_516_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_517_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_517_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_518_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_518_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_519_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_519_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_520_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_520_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_521_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_521_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_en; // @[lib.scala 343:22]
  wire  _T_21 = io_dec_bp_dec_tlu_flush_leak_one_wb & io_dec_tlu_flush_lower_wb; // @[ifu_bp_ctl.scala 135:54]
  reg  leak_one_f_d1; // @[Reg.scala 27:20]
  wire  _T_22 = ~io_dec_tlu_flush_lower_wb; // @[ifu_bp_ctl.scala 135:102]
  wire  _T_23 = leak_one_f_d1 & _T_22; // @[ifu_bp_ctl.scala 135:100]
  wire  leak_one_f = _T_21 | _T_23; // @[ifu_bp_ctl.scala 135:83]
  wire  _T = ~leak_one_f; // @[ifu_bp_ctl.scala 82:58]
  wire  exu_mp_valid = io_exu_bp_exu_mp_pkt_bits_misp & _T; // @[ifu_bp_ctl.scala 82:56]
  wire  dec_tlu_error_wb = io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error | io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu_bp_ctl.scala 105:50]
  wire [7:0] _T_4 = io_ifc_fetch_addr_f[8:1] ^ io_ifc_fetch_addr_f[16:9]; // @[lib.scala 51:47]
  wire [7:0] btb_rd_addr_f = _T_4 ^ io_ifc_fetch_addr_f[24:17]; // @[lib.scala 51:85]
  wire [29:0] fetch_addr_p1_f = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[ifu_bp_ctl.scala 113:51]
  wire [30:0] _T_8 = {fetch_addr_p1_f,1'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_11 = _T_8[8:1] ^ _T_8[16:9]; // @[lib.scala 51:47]
  wire [7:0] btb_rd_addr_p1_f = _T_11 ^ _T_8[24:17]; // @[lib.scala 51:85]
  wire  _T_162 = ~io_ifc_fetch_addr_f[0]; // @[ifu_bp_ctl.scala 191:37]
  wire  _T_2690 = btb_rd_addr_f == 8'h0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_645; // @[Reg.scala 27:20]
  wire [21:0] _T_3202 = _T_2690 ? _T_645 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_2692 = btb_rd_addr_f == 8'h1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_649; // @[Reg.scala 27:20]
  wire [21:0] _T_3203 = _T_2692 ? _T_649 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3458 = _T_3202 | _T_3203; // @[Mux.scala 27:72]
  wire  _T_2694 = btb_rd_addr_f == 8'h2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_653; // @[Reg.scala 27:20]
  wire [21:0] _T_3204 = _T_2694 ? _T_653 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3459 = _T_3458 | _T_3204; // @[Mux.scala 27:72]
  wire  _T_2696 = btb_rd_addr_f == 8'h3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_657; // @[Reg.scala 27:20]
  wire [21:0] _T_3205 = _T_2696 ? _T_657 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3460 = _T_3459 | _T_3205; // @[Mux.scala 27:72]
  wire  _T_2698 = btb_rd_addr_f == 8'h4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_661; // @[Reg.scala 27:20]
  wire [21:0] _T_3206 = _T_2698 ? _T_661 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3461 = _T_3460 | _T_3206; // @[Mux.scala 27:72]
  wire  _T_2700 = btb_rd_addr_f == 8'h5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_665; // @[Reg.scala 27:20]
  wire [21:0] _T_3207 = _T_2700 ? _T_665 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3462 = _T_3461 | _T_3207; // @[Mux.scala 27:72]
  wire  _T_2702 = btb_rd_addr_f == 8'h6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_669; // @[Reg.scala 27:20]
  wire [21:0] _T_3208 = _T_2702 ? _T_669 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3463 = _T_3462 | _T_3208; // @[Mux.scala 27:72]
  wire  _T_2704 = btb_rd_addr_f == 8'h7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_673; // @[Reg.scala 27:20]
  wire [21:0] _T_3209 = _T_2704 ? _T_673 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3464 = _T_3463 | _T_3209; // @[Mux.scala 27:72]
  wire  _T_2706 = btb_rd_addr_f == 8'h8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_677; // @[Reg.scala 27:20]
  wire [21:0] _T_3210 = _T_2706 ? _T_677 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3465 = _T_3464 | _T_3210; // @[Mux.scala 27:72]
  wire  _T_2708 = btb_rd_addr_f == 8'h9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_681; // @[Reg.scala 27:20]
  wire [21:0] _T_3211 = _T_2708 ? _T_681 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3466 = _T_3465 | _T_3211; // @[Mux.scala 27:72]
  wire  _T_2710 = btb_rd_addr_f == 8'ha; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_685; // @[Reg.scala 27:20]
  wire [21:0] _T_3212 = _T_2710 ? _T_685 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3467 = _T_3466 | _T_3212; // @[Mux.scala 27:72]
  wire  _T_2712 = btb_rd_addr_f == 8'hb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_689; // @[Reg.scala 27:20]
  wire [21:0] _T_3213 = _T_2712 ? _T_689 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3468 = _T_3467 | _T_3213; // @[Mux.scala 27:72]
  wire  _T_2714 = btb_rd_addr_f == 8'hc; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_693; // @[Reg.scala 27:20]
  wire [21:0] _T_3214 = _T_2714 ? _T_693 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3469 = _T_3468 | _T_3214; // @[Mux.scala 27:72]
  wire  _T_2716 = btb_rd_addr_f == 8'hd; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_697; // @[Reg.scala 27:20]
  wire [21:0] _T_3215 = _T_2716 ? _T_697 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3470 = _T_3469 | _T_3215; // @[Mux.scala 27:72]
  wire  _T_2718 = btb_rd_addr_f == 8'he; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_701; // @[Reg.scala 27:20]
  wire [21:0] _T_3216 = _T_2718 ? _T_701 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3471 = _T_3470 | _T_3216; // @[Mux.scala 27:72]
  wire  _T_2720 = btb_rd_addr_f == 8'hf; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_705; // @[Reg.scala 27:20]
  wire [21:0] _T_3217 = _T_2720 ? _T_705 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3472 = _T_3471 | _T_3217; // @[Mux.scala 27:72]
  wire  _T_2722 = btb_rd_addr_f == 8'h10; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_709; // @[Reg.scala 27:20]
  wire [21:0] _T_3218 = _T_2722 ? _T_709 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3473 = _T_3472 | _T_3218; // @[Mux.scala 27:72]
  wire  _T_2724 = btb_rd_addr_f == 8'h11; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_713; // @[Reg.scala 27:20]
  wire [21:0] _T_3219 = _T_2724 ? _T_713 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3474 = _T_3473 | _T_3219; // @[Mux.scala 27:72]
  wire  _T_2726 = btb_rd_addr_f == 8'h12; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_717; // @[Reg.scala 27:20]
  wire [21:0] _T_3220 = _T_2726 ? _T_717 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3475 = _T_3474 | _T_3220; // @[Mux.scala 27:72]
  wire  _T_2728 = btb_rd_addr_f == 8'h13; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_721; // @[Reg.scala 27:20]
  wire [21:0] _T_3221 = _T_2728 ? _T_721 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3476 = _T_3475 | _T_3221; // @[Mux.scala 27:72]
  wire  _T_2730 = btb_rd_addr_f == 8'h14; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_725; // @[Reg.scala 27:20]
  wire [21:0] _T_3222 = _T_2730 ? _T_725 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3477 = _T_3476 | _T_3222; // @[Mux.scala 27:72]
  wire  _T_2732 = btb_rd_addr_f == 8'h15; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_729; // @[Reg.scala 27:20]
  wire [21:0] _T_3223 = _T_2732 ? _T_729 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3478 = _T_3477 | _T_3223; // @[Mux.scala 27:72]
  wire  _T_2734 = btb_rd_addr_f == 8'h16; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_733; // @[Reg.scala 27:20]
  wire [21:0] _T_3224 = _T_2734 ? _T_733 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3479 = _T_3478 | _T_3224; // @[Mux.scala 27:72]
  wire  _T_2736 = btb_rd_addr_f == 8'h17; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_737; // @[Reg.scala 27:20]
  wire [21:0] _T_3225 = _T_2736 ? _T_737 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3480 = _T_3479 | _T_3225; // @[Mux.scala 27:72]
  wire  _T_2738 = btb_rd_addr_f == 8'h18; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_741; // @[Reg.scala 27:20]
  wire [21:0] _T_3226 = _T_2738 ? _T_741 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3481 = _T_3480 | _T_3226; // @[Mux.scala 27:72]
  wire  _T_2740 = btb_rd_addr_f == 8'h19; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_745; // @[Reg.scala 27:20]
  wire [21:0] _T_3227 = _T_2740 ? _T_745 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3482 = _T_3481 | _T_3227; // @[Mux.scala 27:72]
  wire  _T_2742 = btb_rd_addr_f == 8'h1a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_749; // @[Reg.scala 27:20]
  wire [21:0] _T_3228 = _T_2742 ? _T_749 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3483 = _T_3482 | _T_3228; // @[Mux.scala 27:72]
  wire  _T_2744 = btb_rd_addr_f == 8'h1b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_753; // @[Reg.scala 27:20]
  wire [21:0] _T_3229 = _T_2744 ? _T_753 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3484 = _T_3483 | _T_3229; // @[Mux.scala 27:72]
  wire  _T_2746 = btb_rd_addr_f == 8'h1c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_757; // @[Reg.scala 27:20]
  wire [21:0] _T_3230 = _T_2746 ? _T_757 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3485 = _T_3484 | _T_3230; // @[Mux.scala 27:72]
  wire  _T_2748 = btb_rd_addr_f == 8'h1d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_761; // @[Reg.scala 27:20]
  wire [21:0] _T_3231 = _T_2748 ? _T_761 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3486 = _T_3485 | _T_3231; // @[Mux.scala 27:72]
  wire  _T_2750 = btb_rd_addr_f == 8'h1e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_765; // @[Reg.scala 27:20]
  wire [21:0] _T_3232 = _T_2750 ? _T_765 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3487 = _T_3486 | _T_3232; // @[Mux.scala 27:72]
  wire  _T_2752 = btb_rd_addr_f == 8'h1f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_769; // @[Reg.scala 27:20]
  wire [21:0] _T_3233 = _T_2752 ? _T_769 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3488 = _T_3487 | _T_3233; // @[Mux.scala 27:72]
  wire  _T_2754 = btb_rd_addr_f == 8'h20; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_773; // @[Reg.scala 27:20]
  wire [21:0] _T_3234 = _T_2754 ? _T_773 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3489 = _T_3488 | _T_3234; // @[Mux.scala 27:72]
  wire  _T_2756 = btb_rd_addr_f == 8'h21; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_777; // @[Reg.scala 27:20]
  wire [21:0] _T_3235 = _T_2756 ? _T_777 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3490 = _T_3489 | _T_3235; // @[Mux.scala 27:72]
  wire  _T_2758 = btb_rd_addr_f == 8'h22; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_781; // @[Reg.scala 27:20]
  wire [21:0] _T_3236 = _T_2758 ? _T_781 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3491 = _T_3490 | _T_3236; // @[Mux.scala 27:72]
  wire  _T_2760 = btb_rd_addr_f == 8'h23; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_785; // @[Reg.scala 27:20]
  wire [21:0] _T_3237 = _T_2760 ? _T_785 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3492 = _T_3491 | _T_3237; // @[Mux.scala 27:72]
  wire  _T_2762 = btb_rd_addr_f == 8'h24; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_789; // @[Reg.scala 27:20]
  wire [21:0] _T_3238 = _T_2762 ? _T_789 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3493 = _T_3492 | _T_3238; // @[Mux.scala 27:72]
  wire  _T_2764 = btb_rd_addr_f == 8'h25; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_793; // @[Reg.scala 27:20]
  wire [21:0] _T_3239 = _T_2764 ? _T_793 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3494 = _T_3493 | _T_3239; // @[Mux.scala 27:72]
  wire  _T_2766 = btb_rd_addr_f == 8'h26; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_797; // @[Reg.scala 27:20]
  wire [21:0] _T_3240 = _T_2766 ? _T_797 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3495 = _T_3494 | _T_3240; // @[Mux.scala 27:72]
  wire  _T_2768 = btb_rd_addr_f == 8'h27; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_801; // @[Reg.scala 27:20]
  wire [21:0] _T_3241 = _T_2768 ? _T_801 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3496 = _T_3495 | _T_3241; // @[Mux.scala 27:72]
  wire  _T_2770 = btb_rd_addr_f == 8'h28; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_805; // @[Reg.scala 27:20]
  wire [21:0] _T_3242 = _T_2770 ? _T_805 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3497 = _T_3496 | _T_3242; // @[Mux.scala 27:72]
  wire  _T_2772 = btb_rd_addr_f == 8'h29; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_809; // @[Reg.scala 27:20]
  wire [21:0] _T_3243 = _T_2772 ? _T_809 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3498 = _T_3497 | _T_3243; // @[Mux.scala 27:72]
  wire  _T_2774 = btb_rd_addr_f == 8'h2a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_813; // @[Reg.scala 27:20]
  wire [21:0] _T_3244 = _T_2774 ? _T_813 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3499 = _T_3498 | _T_3244; // @[Mux.scala 27:72]
  wire  _T_2776 = btb_rd_addr_f == 8'h2b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_817; // @[Reg.scala 27:20]
  wire [21:0] _T_3245 = _T_2776 ? _T_817 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3500 = _T_3499 | _T_3245; // @[Mux.scala 27:72]
  wire  _T_2778 = btb_rd_addr_f == 8'h2c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_821; // @[Reg.scala 27:20]
  wire [21:0] _T_3246 = _T_2778 ? _T_821 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3501 = _T_3500 | _T_3246; // @[Mux.scala 27:72]
  wire  _T_2780 = btb_rd_addr_f == 8'h2d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_825; // @[Reg.scala 27:20]
  wire [21:0] _T_3247 = _T_2780 ? _T_825 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3502 = _T_3501 | _T_3247; // @[Mux.scala 27:72]
  wire  _T_2782 = btb_rd_addr_f == 8'h2e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_829; // @[Reg.scala 27:20]
  wire [21:0] _T_3248 = _T_2782 ? _T_829 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3503 = _T_3502 | _T_3248; // @[Mux.scala 27:72]
  wire  _T_2784 = btb_rd_addr_f == 8'h2f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_833; // @[Reg.scala 27:20]
  wire [21:0] _T_3249 = _T_2784 ? _T_833 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3504 = _T_3503 | _T_3249; // @[Mux.scala 27:72]
  wire  _T_2786 = btb_rd_addr_f == 8'h30; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_837; // @[Reg.scala 27:20]
  wire [21:0] _T_3250 = _T_2786 ? _T_837 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3505 = _T_3504 | _T_3250; // @[Mux.scala 27:72]
  wire  _T_2788 = btb_rd_addr_f == 8'h31; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_841; // @[Reg.scala 27:20]
  wire [21:0] _T_3251 = _T_2788 ? _T_841 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3506 = _T_3505 | _T_3251; // @[Mux.scala 27:72]
  wire  _T_2790 = btb_rd_addr_f == 8'h32; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_845; // @[Reg.scala 27:20]
  wire [21:0] _T_3252 = _T_2790 ? _T_845 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3507 = _T_3506 | _T_3252; // @[Mux.scala 27:72]
  wire  _T_2792 = btb_rd_addr_f == 8'h33; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_849; // @[Reg.scala 27:20]
  wire [21:0] _T_3253 = _T_2792 ? _T_849 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3508 = _T_3507 | _T_3253; // @[Mux.scala 27:72]
  wire  _T_2794 = btb_rd_addr_f == 8'h34; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_853; // @[Reg.scala 27:20]
  wire [21:0] _T_3254 = _T_2794 ? _T_853 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3509 = _T_3508 | _T_3254; // @[Mux.scala 27:72]
  wire  _T_2796 = btb_rd_addr_f == 8'h35; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_857; // @[Reg.scala 27:20]
  wire [21:0] _T_3255 = _T_2796 ? _T_857 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3510 = _T_3509 | _T_3255; // @[Mux.scala 27:72]
  wire  _T_2798 = btb_rd_addr_f == 8'h36; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_861; // @[Reg.scala 27:20]
  wire [21:0] _T_3256 = _T_2798 ? _T_861 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3511 = _T_3510 | _T_3256; // @[Mux.scala 27:72]
  wire  _T_2800 = btb_rd_addr_f == 8'h37; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_865; // @[Reg.scala 27:20]
  wire [21:0] _T_3257 = _T_2800 ? _T_865 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3512 = _T_3511 | _T_3257; // @[Mux.scala 27:72]
  wire  _T_2802 = btb_rd_addr_f == 8'h38; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_869; // @[Reg.scala 27:20]
  wire [21:0] _T_3258 = _T_2802 ? _T_869 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3513 = _T_3512 | _T_3258; // @[Mux.scala 27:72]
  wire  _T_2804 = btb_rd_addr_f == 8'h39; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_873; // @[Reg.scala 27:20]
  wire [21:0] _T_3259 = _T_2804 ? _T_873 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3514 = _T_3513 | _T_3259; // @[Mux.scala 27:72]
  wire  _T_2806 = btb_rd_addr_f == 8'h3a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_877; // @[Reg.scala 27:20]
  wire [21:0] _T_3260 = _T_2806 ? _T_877 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3515 = _T_3514 | _T_3260; // @[Mux.scala 27:72]
  wire  _T_2808 = btb_rd_addr_f == 8'h3b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_881; // @[Reg.scala 27:20]
  wire [21:0] _T_3261 = _T_2808 ? _T_881 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3516 = _T_3515 | _T_3261; // @[Mux.scala 27:72]
  wire  _T_2810 = btb_rd_addr_f == 8'h3c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_885; // @[Reg.scala 27:20]
  wire [21:0] _T_3262 = _T_2810 ? _T_885 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3517 = _T_3516 | _T_3262; // @[Mux.scala 27:72]
  wire  _T_2812 = btb_rd_addr_f == 8'h3d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_889; // @[Reg.scala 27:20]
  wire [21:0] _T_3263 = _T_2812 ? _T_889 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3518 = _T_3517 | _T_3263; // @[Mux.scala 27:72]
  wire  _T_2814 = btb_rd_addr_f == 8'h3e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_893; // @[Reg.scala 27:20]
  wire [21:0] _T_3264 = _T_2814 ? _T_893 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3519 = _T_3518 | _T_3264; // @[Mux.scala 27:72]
  wire  _T_2816 = btb_rd_addr_f == 8'h3f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_897; // @[Reg.scala 27:20]
  wire [21:0] _T_3265 = _T_2816 ? _T_897 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3520 = _T_3519 | _T_3265; // @[Mux.scala 27:72]
  wire  _T_2818 = btb_rd_addr_f == 8'h40; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_901; // @[Reg.scala 27:20]
  wire [21:0] _T_3266 = _T_2818 ? _T_901 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3521 = _T_3520 | _T_3266; // @[Mux.scala 27:72]
  wire  _T_2820 = btb_rd_addr_f == 8'h41; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_905; // @[Reg.scala 27:20]
  wire [21:0] _T_3267 = _T_2820 ? _T_905 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3522 = _T_3521 | _T_3267; // @[Mux.scala 27:72]
  wire  _T_2822 = btb_rd_addr_f == 8'h42; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_909; // @[Reg.scala 27:20]
  wire [21:0] _T_3268 = _T_2822 ? _T_909 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3523 = _T_3522 | _T_3268; // @[Mux.scala 27:72]
  wire  _T_2824 = btb_rd_addr_f == 8'h43; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_913; // @[Reg.scala 27:20]
  wire [21:0] _T_3269 = _T_2824 ? _T_913 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3524 = _T_3523 | _T_3269; // @[Mux.scala 27:72]
  wire  _T_2826 = btb_rd_addr_f == 8'h44; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_917; // @[Reg.scala 27:20]
  wire [21:0] _T_3270 = _T_2826 ? _T_917 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3525 = _T_3524 | _T_3270; // @[Mux.scala 27:72]
  wire  _T_2828 = btb_rd_addr_f == 8'h45; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_921; // @[Reg.scala 27:20]
  wire [21:0] _T_3271 = _T_2828 ? _T_921 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3526 = _T_3525 | _T_3271; // @[Mux.scala 27:72]
  wire  _T_2830 = btb_rd_addr_f == 8'h46; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_925; // @[Reg.scala 27:20]
  wire [21:0] _T_3272 = _T_2830 ? _T_925 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3527 = _T_3526 | _T_3272; // @[Mux.scala 27:72]
  wire  _T_2832 = btb_rd_addr_f == 8'h47; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_929; // @[Reg.scala 27:20]
  wire [21:0] _T_3273 = _T_2832 ? _T_929 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3528 = _T_3527 | _T_3273; // @[Mux.scala 27:72]
  wire  _T_2834 = btb_rd_addr_f == 8'h48; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_933; // @[Reg.scala 27:20]
  wire [21:0] _T_3274 = _T_2834 ? _T_933 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3529 = _T_3528 | _T_3274; // @[Mux.scala 27:72]
  wire  _T_2836 = btb_rd_addr_f == 8'h49; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_937; // @[Reg.scala 27:20]
  wire [21:0] _T_3275 = _T_2836 ? _T_937 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3530 = _T_3529 | _T_3275; // @[Mux.scala 27:72]
  wire  _T_2838 = btb_rd_addr_f == 8'h4a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_941; // @[Reg.scala 27:20]
  wire [21:0] _T_3276 = _T_2838 ? _T_941 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3531 = _T_3530 | _T_3276; // @[Mux.scala 27:72]
  wire  _T_2840 = btb_rd_addr_f == 8'h4b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_945; // @[Reg.scala 27:20]
  wire [21:0] _T_3277 = _T_2840 ? _T_945 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3532 = _T_3531 | _T_3277; // @[Mux.scala 27:72]
  wire  _T_2842 = btb_rd_addr_f == 8'h4c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_949; // @[Reg.scala 27:20]
  wire [21:0] _T_3278 = _T_2842 ? _T_949 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3533 = _T_3532 | _T_3278; // @[Mux.scala 27:72]
  wire  _T_2844 = btb_rd_addr_f == 8'h4d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_953; // @[Reg.scala 27:20]
  wire [21:0] _T_3279 = _T_2844 ? _T_953 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3534 = _T_3533 | _T_3279; // @[Mux.scala 27:72]
  wire  _T_2846 = btb_rd_addr_f == 8'h4e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_957; // @[Reg.scala 27:20]
  wire [21:0] _T_3280 = _T_2846 ? _T_957 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3535 = _T_3534 | _T_3280; // @[Mux.scala 27:72]
  wire  _T_2848 = btb_rd_addr_f == 8'h4f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_961; // @[Reg.scala 27:20]
  wire [21:0] _T_3281 = _T_2848 ? _T_961 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3536 = _T_3535 | _T_3281; // @[Mux.scala 27:72]
  wire  _T_2850 = btb_rd_addr_f == 8'h50; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_965; // @[Reg.scala 27:20]
  wire [21:0] _T_3282 = _T_2850 ? _T_965 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3537 = _T_3536 | _T_3282; // @[Mux.scala 27:72]
  wire  _T_2852 = btb_rd_addr_f == 8'h51; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_969; // @[Reg.scala 27:20]
  wire [21:0] _T_3283 = _T_2852 ? _T_969 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3538 = _T_3537 | _T_3283; // @[Mux.scala 27:72]
  wire  _T_2854 = btb_rd_addr_f == 8'h52; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_973; // @[Reg.scala 27:20]
  wire [21:0] _T_3284 = _T_2854 ? _T_973 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3539 = _T_3538 | _T_3284; // @[Mux.scala 27:72]
  wire  _T_2856 = btb_rd_addr_f == 8'h53; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_977; // @[Reg.scala 27:20]
  wire [21:0] _T_3285 = _T_2856 ? _T_977 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3540 = _T_3539 | _T_3285; // @[Mux.scala 27:72]
  wire  _T_2858 = btb_rd_addr_f == 8'h54; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_981; // @[Reg.scala 27:20]
  wire [21:0] _T_3286 = _T_2858 ? _T_981 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3541 = _T_3540 | _T_3286; // @[Mux.scala 27:72]
  wire  _T_2860 = btb_rd_addr_f == 8'h55; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_985; // @[Reg.scala 27:20]
  wire [21:0] _T_3287 = _T_2860 ? _T_985 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3542 = _T_3541 | _T_3287; // @[Mux.scala 27:72]
  wire  _T_2862 = btb_rd_addr_f == 8'h56; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_989; // @[Reg.scala 27:20]
  wire [21:0] _T_3288 = _T_2862 ? _T_989 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3543 = _T_3542 | _T_3288; // @[Mux.scala 27:72]
  wire  _T_2864 = btb_rd_addr_f == 8'h57; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_993; // @[Reg.scala 27:20]
  wire [21:0] _T_3289 = _T_2864 ? _T_993 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3544 = _T_3543 | _T_3289; // @[Mux.scala 27:72]
  wire  _T_2866 = btb_rd_addr_f == 8'h58; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_997; // @[Reg.scala 27:20]
  wire [21:0] _T_3290 = _T_2866 ? _T_997 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3545 = _T_3544 | _T_3290; // @[Mux.scala 27:72]
  wire  _T_2868 = btb_rd_addr_f == 8'h59; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1001; // @[Reg.scala 27:20]
  wire [21:0] _T_3291 = _T_2868 ? _T_1001 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3546 = _T_3545 | _T_3291; // @[Mux.scala 27:72]
  wire  _T_2870 = btb_rd_addr_f == 8'h5a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1005; // @[Reg.scala 27:20]
  wire [21:0] _T_3292 = _T_2870 ? _T_1005 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3547 = _T_3546 | _T_3292; // @[Mux.scala 27:72]
  wire  _T_2872 = btb_rd_addr_f == 8'h5b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1009; // @[Reg.scala 27:20]
  wire [21:0] _T_3293 = _T_2872 ? _T_1009 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3548 = _T_3547 | _T_3293; // @[Mux.scala 27:72]
  wire  _T_2874 = btb_rd_addr_f == 8'h5c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1013; // @[Reg.scala 27:20]
  wire [21:0] _T_3294 = _T_2874 ? _T_1013 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3549 = _T_3548 | _T_3294; // @[Mux.scala 27:72]
  wire  _T_2876 = btb_rd_addr_f == 8'h5d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1017; // @[Reg.scala 27:20]
  wire [21:0] _T_3295 = _T_2876 ? _T_1017 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3550 = _T_3549 | _T_3295; // @[Mux.scala 27:72]
  wire  _T_2878 = btb_rd_addr_f == 8'h5e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1021; // @[Reg.scala 27:20]
  wire [21:0] _T_3296 = _T_2878 ? _T_1021 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3551 = _T_3550 | _T_3296; // @[Mux.scala 27:72]
  wire  _T_2880 = btb_rd_addr_f == 8'h5f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1025; // @[Reg.scala 27:20]
  wire [21:0] _T_3297 = _T_2880 ? _T_1025 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3552 = _T_3551 | _T_3297; // @[Mux.scala 27:72]
  wire  _T_2882 = btb_rd_addr_f == 8'h60; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1029; // @[Reg.scala 27:20]
  wire [21:0] _T_3298 = _T_2882 ? _T_1029 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3553 = _T_3552 | _T_3298; // @[Mux.scala 27:72]
  wire  _T_2884 = btb_rd_addr_f == 8'h61; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1033; // @[Reg.scala 27:20]
  wire [21:0] _T_3299 = _T_2884 ? _T_1033 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3554 = _T_3553 | _T_3299; // @[Mux.scala 27:72]
  wire  _T_2886 = btb_rd_addr_f == 8'h62; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1037; // @[Reg.scala 27:20]
  wire [21:0] _T_3300 = _T_2886 ? _T_1037 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3555 = _T_3554 | _T_3300; // @[Mux.scala 27:72]
  wire  _T_2888 = btb_rd_addr_f == 8'h63; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1041; // @[Reg.scala 27:20]
  wire [21:0] _T_3301 = _T_2888 ? _T_1041 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3556 = _T_3555 | _T_3301; // @[Mux.scala 27:72]
  wire  _T_2890 = btb_rd_addr_f == 8'h64; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1045; // @[Reg.scala 27:20]
  wire [21:0] _T_3302 = _T_2890 ? _T_1045 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3557 = _T_3556 | _T_3302; // @[Mux.scala 27:72]
  wire  _T_2892 = btb_rd_addr_f == 8'h65; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1049; // @[Reg.scala 27:20]
  wire [21:0] _T_3303 = _T_2892 ? _T_1049 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3558 = _T_3557 | _T_3303; // @[Mux.scala 27:72]
  wire  _T_2894 = btb_rd_addr_f == 8'h66; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1053; // @[Reg.scala 27:20]
  wire [21:0] _T_3304 = _T_2894 ? _T_1053 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3559 = _T_3558 | _T_3304; // @[Mux.scala 27:72]
  wire  _T_2896 = btb_rd_addr_f == 8'h67; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1057; // @[Reg.scala 27:20]
  wire [21:0] _T_3305 = _T_2896 ? _T_1057 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3560 = _T_3559 | _T_3305; // @[Mux.scala 27:72]
  wire  _T_2898 = btb_rd_addr_f == 8'h68; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1061; // @[Reg.scala 27:20]
  wire [21:0] _T_3306 = _T_2898 ? _T_1061 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3561 = _T_3560 | _T_3306; // @[Mux.scala 27:72]
  wire  _T_2900 = btb_rd_addr_f == 8'h69; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1065; // @[Reg.scala 27:20]
  wire [21:0] _T_3307 = _T_2900 ? _T_1065 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3562 = _T_3561 | _T_3307; // @[Mux.scala 27:72]
  wire  _T_2902 = btb_rd_addr_f == 8'h6a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1069; // @[Reg.scala 27:20]
  wire [21:0] _T_3308 = _T_2902 ? _T_1069 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3563 = _T_3562 | _T_3308; // @[Mux.scala 27:72]
  wire  _T_2904 = btb_rd_addr_f == 8'h6b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1073; // @[Reg.scala 27:20]
  wire [21:0] _T_3309 = _T_2904 ? _T_1073 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3564 = _T_3563 | _T_3309; // @[Mux.scala 27:72]
  wire  _T_2906 = btb_rd_addr_f == 8'h6c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1077; // @[Reg.scala 27:20]
  wire [21:0] _T_3310 = _T_2906 ? _T_1077 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3565 = _T_3564 | _T_3310; // @[Mux.scala 27:72]
  wire  _T_2908 = btb_rd_addr_f == 8'h6d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1081; // @[Reg.scala 27:20]
  wire [21:0] _T_3311 = _T_2908 ? _T_1081 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3566 = _T_3565 | _T_3311; // @[Mux.scala 27:72]
  wire  _T_2910 = btb_rd_addr_f == 8'h6e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1085; // @[Reg.scala 27:20]
  wire [21:0] _T_3312 = _T_2910 ? _T_1085 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3567 = _T_3566 | _T_3312; // @[Mux.scala 27:72]
  wire  _T_2912 = btb_rd_addr_f == 8'h6f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1089; // @[Reg.scala 27:20]
  wire [21:0] _T_3313 = _T_2912 ? _T_1089 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3568 = _T_3567 | _T_3313; // @[Mux.scala 27:72]
  wire  _T_2914 = btb_rd_addr_f == 8'h70; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1093; // @[Reg.scala 27:20]
  wire [21:0] _T_3314 = _T_2914 ? _T_1093 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3569 = _T_3568 | _T_3314; // @[Mux.scala 27:72]
  wire  _T_2916 = btb_rd_addr_f == 8'h71; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1097; // @[Reg.scala 27:20]
  wire [21:0] _T_3315 = _T_2916 ? _T_1097 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3570 = _T_3569 | _T_3315; // @[Mux.scala 27:72]
  wire  _T_2918 = btb_rd_addr_f == 8'h72; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1101; // @[Reg.scala 27:20]
  wire [21:0] _T_3316 = _T_2918 ? _T_1101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3571 = _T_3570 | _T_3316; // @[Mux.scala 27:72]
  wire  _T_2920 = btb_rd_addr_f == 8'h73; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1105; // @[Reg.scala 27:20]
  wire [21:0] _T_3317 = _T_2920 ? _T_1105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3572 = _T_3571 | _T_3317; // @[Mux.scala 27:72]
  wire  _T_2922 = btb_rd_addr_f == 8'h74; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1109; // @[Reg.scala 27:20]
  wire [21:0] _T_3318 = _T_2922 ? _T_1109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3573 = _T_3572 | _T_3318; // @[Mux.scala 27:72]
  wire  _T_2924 = btb_rd_addr_f == 8'h75; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1113; // @[Reg.scala 27:20]
  wire [21:0] _T_3319 = _T_2924 ? _T_1113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3574 = _T_3573 | _T_3319; // @[Mux.scala 27:72]
  wire  _T_2926 = btb_rd_addr_f == 8'h76; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1117; // @[Reg.scala 27:20]
  wire [21:0] _T_3320 = _T_2926 ? _T_1117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3575 = _T_3574 | _T_3320; // @[Mux.scala 27:72]
  wire  _T_2928 = btb_rd_addr_f == 8'h77; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1121; // @[Reg.scala 27:20]
  wire [21:0] _T_3321 = _T_2928 ? _T_1121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3576 = _T_3575 | _T_3321; // @[Mux.scala 27:72]
  wire  _T_2930 = btb_rd_addr_f == 8'h78; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1125; // @[Reg.scala 27:20]
  wire [21:0] _T_3322 = _T_2930 ? _T_1125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3577 = _T_3576 | _T_3322; // @[Mux.scala 27:72]
  wire  _T_2932 = btb_rd_addr_f == 8'h79; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1129; // @[Reg.scala 27:20]
  wire [21:0] _T_3323 = _T_2932 ? _T_1129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3578 = _T_3577 | _T_3323; // @[Mux.scala 27:72]
  wire  _T_2934 = btb_rd_addr_f == 8'h7a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1133; // @[Reg.scala 27:20]
  wire [21:0] _T_3324 = _T_2934 ? _T_1133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3579 = _T_3578 | _T_3324; // @[Mux.scala 27:72]
  wire  _T_2936 = btb_rd_addr_f == 8'h7b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1137; // @[Reg.scala 27:20]
  wire [21:0] _T_3325 = _T_2936 ? _T_1137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3580 = _T_3579 | _T_3325; // @[Mux.scala 27:72]
  wire  _T_2938 = btb_rd_addr_f == 8'h7c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1141; // @[Reg.scala 27:20]
  wire [21:0] _T_3326 = _T_2938 ? _T_1141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3581 = _T_3580 | _T_3326; // @[Mux.scala 27:72]
  wire  _T_2940 = btb_rd_addr_f == 8'h7d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1145; // @[Reg.scala 27:20]
  wire [21:0] _T_3327 = _T_2940 ? _T_1145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3582 = _T_3581 | _T_3327; // @[Mux.scala 27:72]
  wire  _T_2942 = btb_rd_addr_f == 8'h7e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1149; // @[Reg.scala 27:20]
  wire [21:0] _T_3328 = _T_2942 ? _T_1149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3583 = _T_3582 | _T_3328; // @[Mux.scala 27:72]
  wire  _T_2944 = btb_rd_addr_f == 8'h7f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1153; // @[Reg.scala 27:20]
  wire [21:0] _T_3329 = _T_2944 ? _T_1153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3584 = _T_3583 | _T_3329; // @[Mux.scala 27:72]
  wire  _T_2946 = btb_rd_addr_f == 8'h80; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1157; // @[Reg.scala 27:20]
  wire [21:0] _T_3330 = _T_2946 ? _T_1157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3585 = _T_3584 | _T_3330; // @[Mux.scala 27:72]
  wire  _T_2948 = btb_rd_addr_f == 8'h81; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1161; // @[Reg.scala 27:20]
  wire [21:0] _T_3331 = _T_2948 ? _T_1161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3586 = _T_3585 | _T_3331; // @[Mux.scala 27:72]
  wire  _T_2950 = btb_rd_addr_f == 8'h82; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1165; // @[Reg.scala 27:20]
  wire [21:0] _T_3332 = _T_2950 ? _T_1165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3587 = _T_3586 | _T_3332; // @[Mux.scala 27:72]
  wire  _T_2952 = btb_rd_addr_f == 8'h83; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1169; // @[Reg.scala 27:20]
  wire [21:0] _T_3333 = _T_2952 ? _T_1169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3588 = _T_3587 | _T_3333; // @[Mux.scala 27:72]
  wire  _T_2954 = btb_rd_addr_f == 8'h84; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1173; // @[Reg.scala 27:20]
  wire [21:0] _T_3334 = _T_2954 ? _T_1173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3589 = _T_3588 | _T_3334; // @[Mux.scala 27:72]
  wire  _T_2956 = btb_rd_addr_f == 8'h85; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1177; // @[Reg.scala 27:20]
  wire [21:0] _T_3335 = _T_2956 ? _T_1177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3590 = _T_3589 | _T_3335; // @[Mux.scala 27:72]
  wire  _T_2958 = btb_rd_addr_f == 8'h86; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1181; // @[Reg.scala 27:20]
  wire [21:0] _T_3336 = _T_2958 ? _T_1181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3591 = _T_3590 | _T_3336; // @[Mux.scala 27:72]
  wire  _T_2960 = btb_rd_addr_f == 8'h87; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1185; // @[Reg.scala 27:20]
  wire [21:0] _T_3337 = _T_2960 ? _T_1185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3592 = _T_3591 | _T_3337; // @[Mux.scala 27:72]
  wire  _T_2962 = btb_rd_addr_f == 8'h88; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1189; // @[Reg.scala 27:20]
  wire [21:0] _T_3338 = _T_2962 ? _T_1189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3593 = _T_3592 | _T_3338; // @[Mux.scala 27:72]
  wire  _T_2964 = btb_rd_addr_f == 8'h89; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1193; // @[Reg.scala 27:20]
  wire [21:0] _T_3339 = _T_2964 ? _T_1193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3594 = _T_3593 | _T_3339; // @[Mux.scala 27:72]
  wire  _T_2966 = btb_rd_addr_f == 8'h8a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1197; // @[Reg.scala 27:20]
  wire [21:0] _T_3340 = _T_2966 ? _T_1197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3595 = _T_3594 | _T_3340; // @[Mux.scala 27:72]
  wire  _T_2968 = btb_rd_addr_f == 8'h8b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1201; // @[Reg.scala 27:20]
  wire [21:0] _T_3341 = _T_2968 ? _T_1201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3596 = _T_3595 | _T_3341; // @[Mux.scala 27:72]
  wire  _T_2970 = btb_rd_addr_f == 8'h8c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1205; // @[Reg.scala 27:20]
  wire [21:0] _T_3342 = _T_2970 ? _T_1205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3597 = _T_3596 | _T_3342; // @[Mux.scala 27:72]
  wire  _T_2972 = btb_rd_addr_f == 8'h8d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1209; // @[Reg.scala 27:20]
  wire [21:0] _T_3343 = _T_2972 ? _T_1209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3598 = _T_3597 | _T_3343; // @[Mux.scala 27:72]
  wire  _T_2974 = btb_rd_addr_f == 8'h8e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1213; // @[Reg.scala 27:20]
  wire [21:0] _T_3344 = _T_2974 ? _T_1213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3599 = _T_3598 | _T_3344; // @[Mux.scala 27:72]
  wire  _T_2976 = btb_rd_addr_f == 8'h8f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1217; // @[Reg.scala 27:20]
  wire [21:0] _T_3345 = _T_2976 ? _T_1217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3600 = _T_3599 | _T_3345; // @[Mux.scala 27:72]
  wire  _T_2978 = btb_rd_addr_f == 8'h90; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1221; // @[Reg.scala 27:20]
  wire [21:0] _T_3346 = _T_2978 ? _T_1221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3601 = _T_3600 | _T_3346; // @[Mux.scala 27:72]
  wire  _T_2980 = btb_rd_addr_f == 8'h91; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1225; // @[Reg.scala 27:20]
  wire [21:0] _T_3347 = _T_2980 ? _T_1225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3602 = _T_3601 | _T_3347; // @[Mux.scala 27:72]
  wire  _T_2982 = btb_rd_addr_f == 8'h92; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1229; // @[Reg.scala 27:20]
  wire [21:0] _T_3348 = _T_2982 ? _T_1229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3603 = _T_3602 | _T_3348; // @[Mux.scala 27:72]
  wire  _T_2984 = btb_rd_addr_f == 8'h93; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1233; // @[Reg.scala 27:20]
  wire [21:0] _T_3349 = _T_2984 ? _T_1233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3604 = _T_3603 | _T_3349; // @[Mux.scala 27:72]
  wire  _T_2986 = btb_rd_addr_f == 8'h94; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1237; // @[Reg.scala 27:20]
  wire [21:0] _T_3350 = _T_2986 ? _T_1237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3605 = _T_3604 | _T_3350; // @[Mux.scala 27:72]
  wire  _T_2988 = btb_rd_addr_f == 8'h95; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1241; // @[Reg.scala 27:20]
  wire [21:0] _T_3351 = _T_2988 ? _T_1241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3606 = _T_3605 | _T_3351; // @[Mux.scala 27:72]
  wire  _T_2990 = btb_rd_addr_f == 8'h96; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1245; // @[Reg.scala 27:20]
  wire [21:0] _T_3352 = _T_2990 ? _T_1245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3607 = _T_3606 | _T_3352; // @[Mux.scala 27:72]
  wire  _T_2992 = btb_rd_addr_f == 8'h97; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1249; // @[Reg.scala 27:20]
  wire [21:0] _T_3353 = _T_2992 ? _T_1249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3608 = _T_3607 | _T_3353; // @[Mux.scala 27:72]
  wire  _T_2994 = btb_rd_addr_f == 8'h98; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1253; // @[Reg.scala 27:20]
  wire [21:0] _T_3354 = _T_2994 ? _T_1253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3609 = _T_3608 | _T_3354; // @[Mux.scala 27:72]
  wire  _T_2996 = btb_rd_addr_f == 8'h99; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1257; // @[Reg.scala 27:20]
  wire [21:0] _T_3355 = _T_2996 ? _T_1257 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3610 = _T_3609 | _T_3355; // @[Mux.scala 27:72]
  wire  _T_2998 = btb_rd_addr_f == 8'h9a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1261; // @[Reg.scala 27:20]
  wire [21:0] _T_3356 = _T_2998 ? _T_1261 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3611 = _T_3610 | _T_3356; // @[Mux.scala 27:72]
  wire  _T_3000 = btb_rd_addr_f == 8'h9b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1265; // @[Reg.scala 27:20]
  wire [21:0] _T_3357 = _T_3000 ? _T_1265 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3612 = _T_3611 | _T_3357; // @[Mux.scala 27:72]
  wire  _T_3002 = btb_rd_addr_f == 8'h9c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1269; // @[Reg.scala 27:20]
  wire [21:0] _T_3358 = _T_3002 ? _T_1269 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3613 = _T_3612 | _T_3358; // @[Mux.scala 27:72]
  wire  _T_3004 = btb_rd_addr_f == 8'h9d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1273; // @[Reg.scala 27:20]
  wire [21:0] _T_3359 = _T_3004 ? _T_1273 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3614 = _T_3613 | _T_3359; // @[Mux.scala 27:72]
  wire  _T_3006 = btb_rd_addr_f == 8'h9e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1277; // @[Reg.scala 27:20]
  wire [21:0] _T_3360 = _T_3006 ? _T_1277 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3615 = _T_3614 | _T_3360; // @[Mux.scala 27:72]
  wire  _T_3008 = btb_rd_addr_f == 8'h9f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1281; // @[Reg.scala 27:20]
  wire [21:0] _T_3361 = _T_3008 ? _T_1281 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3616 = _T_3615 | _T_3361; // @[Mux.scala 27:72]
  wire  _T_3010 = btb_rd_addr_f == 8'ha0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1285; // @[Reg.scala 27:20]
  wire [21:0] _T_3362 = _T_3010 ? _T_1285 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3617 = _T_3616 | _T_3362; // @[Mux.scala 27:72]
  wire  _T_3012 = btb_rd_addr_f == 8'ha1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1289; // @[Reg.scala 27:20]
  wire [21:0] _T_3363 = _T_3012 ? _T_1289 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3618 = _T_3617 | _T_3363; // @[Mux.scala 27:72]
  wire  _T_3014 = btb_rd_addr_f == 8'ha2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1293; // @[Reg.scala 27:20]
  wire [21:0] _T_3364 = _T_3014 ? _T_1293 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3619 = _T_3618 | _T_3364; // @[Mux.scala 27:72]
  wire  _T_3016 = btb_rd_addr_f == 8'ha3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1297; // @[Reg.scala 27:20]
  wire [21:0] _T_3365 = _T_3016 ? _T_1297 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3620 = _T_3619 | _T_3365; // @[Mux.scala 27:72]
  wire  _T_3018 = btb_rd_addr_f == 8'ha4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1301; // @[Reg.scala 27:20]
  wire [21:0] _T_3366 = _T_3018 ? _T_1301 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3621 = _T_3620 | _T_3366; // @[Mux.scala 27:72]
  wire  _T_3020 = btb_rd_addr_f == 8'ha5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1305; // @[Reg.scala 27:20]
  wire [21:0] _T_3367 = _T_3020 ? _T_1305 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3622 = _T_3621 | _T_3367; // @[Mux.scala 27:72]
  wire  _T_3022 = btb_rd_addr_f == 8'ha6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1309; // @[Reg.scala 27:20]
  wire [21:0] _T_3368 = _T_3022 ? _T_1309 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3623 = _T_3622 | _T_3368; // @[Mux.scala 27:72]
  wire  _T_3024 = btb_rd_addr_f == 8'ha7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1313; // @[Reg.scala 27:20]
  wire [21:0] _T_3369 = _T_3024 ? _T_1313 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3624 = _T_3623 | _T_3369; // @[Mux.scala 27:72]
  wire  _T_3026 = btb_rd_addr_f == 8'ha8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1317; // @[Reg.scala 27:20]
  wire [21:0] _T_3370 = _T_3026 ? _T_1317 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3625 = _T_3624 | _T_3370; // @[Mux.scala 27:72]
  wire  _T_3028 = btb_rd_addr_f == 8'ha9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1321; // @[Reg.scala 27:20]
  wire [21:0] _T_3371 = _T_3028 ? _T_1321 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3626 = _T_3625 | _T_3371; // @[Mux.scala 27:72]
  wire  _T_3030 = btb_rd_addr_f == 8'haa; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1325; // @[Reg.scala 27:20]
  wire [21:0] _T_3372 = _T_3030 ? _T_1325 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3627 = _T_3626 | _T_3372; // @[Mux.scala 27:72]
  wire  _T_3032 = btb_rd_addr_f == 8'hab; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1329; // @[Reg.scala 27:20]
  wire [21:0] _T_3373 = _T_3032 ? _T_1329 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3628 = _T_3627 | _T_3373; // @[Mux.scala 27:72]
  wire  _T_3034 = btb_rd_addr_f == 8'hac; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1333; // @[Reg.scala 27:20]
  wire [21:0] _T_3374 = _T_3034 ? _T_1333 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3629 = _T_3628 | _T_3374; // @[Mux.scala 27:72]
  wire  _T_3036 = btb_rd_addr_f == 8'had; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1337; // @[Reg.scala 27:20]
  wire [21:0] _T_3375 = _T_3036 ? _T_1337 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3630 = _T_3629 | _T_3375; // @[Mux.scala 27:72]
  wire  _T_3038 = btb_rd_addr_f == 8'hae; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1341; // @[Reg.scala 27:20]
  wire [21:0] _T_3376 = _T_3038 ? _T_1341 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3631 = _T_3630 | _T_3376; // @[Mux.scala 27:72]
  wire  _T_3040 = btb_rd_addr_f == 8'haf; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1345; // @[Reg.scala 27:20]
  wire [21:0] _T_3377 = _T_3040 ? _T_1345 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3632 = _T_3631 | _T_3377; // @[Mux.scala 27:72]
  wire  _T_3042 = btb_rd_addr_f == 8'hb0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1349; // @[Reg.scala 27:20]
  wire [21:0] _T_3378 = _T_3042 ? _T_1349 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3633 = _T_3632 | _T_3378; // @[Mux.scala 27:72]
  wire  _T_3044 = btb_rd_addr_f == 8'hb1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1353; // @[Reg.scala 27:20]
  wire [21:0] _T_3379 = _T_3044 ? _T_1353 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3634 = _T_3633 | _T_3379; // @[Mux.scala 27:72]
  wire  _T_3046 = btb_rd_addr_f == 8'hb2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1357; // @[Reg.scala 27:20]
  wire [21:0] _T_3380 = _T_3046 ? _T_1357 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3635 = _T_3634 | _T_3380; // @[Mux.scala 27:72]
  wire  _T_3048 = btb_rd_addr_f == 8'hb3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1361; // @[Reg.scala 27:20]
  wire [21:0] _T_3381 = _T_3048 ? _T_1361 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3636 = _T_3635 | _T_3381; // @[Mux.scala 27:72]
  wire  _T_3050 = btb_rd_addr_f == 8'hb4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1365; // @[Reg.scala 27:20]
  wire [21:0] _T_3382 = _T_3050 ? _T_1365 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3637 = _T_3636 | _T_3382; // @[Mux.scala 27:72]
  wire  _T_3052 = btb_rd_addr_f == 8'hb5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1369; // @[Reg.scala 27:20]
  wire [21:0] _T_3383 = _T_3052 ? _T_1369 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3638 = _T_3637 | _T_3383; // @[Mux.scala 27:72]
  wire  _T_3054 = btb_rd_addr_f == 8'hb6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1373; // @[Reg.scala 27:20]
  wire [21:0] _T_3384 = _T_3054 ? _T_1373 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3639 = _T_3638 | _T_3384; // @[Mux.scala 27:72]
  wire  _T_3056 = btb_rd_addr_f == 8'hb7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1377; // @[Reg.scala 27:20]
  wire [21:0] _T_3385 = _T_3056 ? _T_1377 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3640 = _T_3639 | _T_3385; // @[Mux.scala 27:72]
  wire  _T_3058 = btb_rd_addr_f == 8'hb8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1381; // @[Reg.scala 27:20]
  wire [21:0] _T_3386 = _T_3058 ? _T_1381 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3641 = _T_3640 | _T_3386; // @[Mux.scala 27:72]
  wire  _T_3060 = btb_rd_addr_f == 8'hb9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1385; // @[Reg.scala 27:20]
  wire [21:0] _T_3387 = _T_3060 ? _T_1385 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3642 = _T_3641 | _T_3387; // @[Mux.scala 27:72]
  wire  _T_3062 = btb_rd_addr_f == 8'hba; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1389; // @[Reg.scala 27:20]
  wire [21:0] _T_3388 = _T_3062 ? _T_1389 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3643 = _T_3642 | _T_3388; // @[Mux.scala 27:72]
  wire  _T_3064 = btb_rd_addr_f == 8'hbb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1393; // @[Reg.scala 27:20]
  wire [21:0] _T_3389 = _T_3064 ? _T_1393 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3644 = _T_3643 | _T_3389; // @[Mux.scala 27:72]
  wire  _T_3066 = btb_rd_addr_f == 8'hbc; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1397; // @[Reg.scala 27:20]
  wire [21:0] _T_3390 = _T_3066 ? _T_1397 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3645 = _T_3644 | _T_3390; // @[Mux.scala 27:72]
  wire  _T_3068 = btb_rd_addr_f == 8'hbd; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1401; // @[Reg.scala 27:20]
  wire [21:0] _T_3391 = _T_3068 ? _T_1401 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3646 = _T_3645 | _T_3391; // @[Mux.scala 27:72]
  wire  _T_3070 = btb_rd_addr_f == 8'hbe; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1405; // @[Reg.scala 27:20]
  wire [21:0] _T_3392 = _T_3070 ? _T_1405 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3647 = _T_3646 | _T_3392; // @[Mux.scala 27:72]
  wire  _T_3072 = btb_rd_addr_f == 8'hbf; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1409; // @[Reg.scala 27:20]
  wire [21:0] _T_3393 = _T_3072 ? _T_1409 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3648 = _T_3647 | _T_3393; // @[Mux.scala 27:72]
  wire  _T_3074 = btb_rd_addr_f == 8'hc0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1413; // @[Reg.scala 27:20]
  wire [21:0] _T_3394 = _T_3074 ? _T_1413 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3649 = _T_3648 | _T_3394; // @[Mux.scala 27:72]
  wire  _T_3076 = btb_rd_addr_f == 8'hc1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1417; // @[Reg.scala 27:20]
  wire [21:0] _T_3395 = _T_3076 ? _T_1417 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3650 = _T_3649 | _T_3395; // @[Mux.scala 27:72]
  wire  _T_3078 = btb_rd_addr_f == 8'hc2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1421; // @[Reg.scala 27:20]
  wire [21:0] _T_3396 = _T_3078 ? _T_1421 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3651 = _T_3650 | _T_3396; // @[Mux.scala 27:72]
  wire  _T_3080 = btb_rd_addr_f == 8'hc3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1425; // @[Reg.scala 27:20]
  wire [21:0] _T_3397 = _T_3080 ? _T_1425 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3652 = _T_3651 | _T_3397; // @[Mux.scala 27:72]
  wire  _T_3082 = btb_rd_addr_f == 8'hc4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1429; // @[Reg.scala 27:20]
  wire [21:0] _T_3398 = _T_3082 ? _T_1429 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3653 = _T_3652 | _T_3398; // @[Mux.scala 27:72]
  wire  _T_3084 = btb_rd_addr_f == 8'hc5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1433; // @[Reg.scala 27:20]
  wire [21:0] _T_3399 = _T_3084 ? _T_1433 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3654 = _T_3653 | _T_3399; // @[Mux.scala 27:72]
  wire  _T_3086 = btb_rd_addr_f == 8'hc6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1437; // @[Reg.scala 27:20]
  wire [21:0] _T_3400 = _T_3086 ? _T_1437 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3655 = _T_3654 | _T_3400; // @[Mux.scala 27:72]
  wire  _T_3088 = btb_rd_addr_f == 8'hc7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1441; // @[Reg.scala 27:20]
  wire [21:0] _T_3401 = _T_3088 ? _T_1441 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3656 = _T_3655 | _T_3401; // @[Mux.scala 27:72]
  wire  _T_3090 = btb_rd_addr_f == 8'hc8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1445; // @[Reg.scala 27:20]
  wire [21:0] _T_3402 = _T_3090 ? _T_1445 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3657 = _T_3656 | _T_3402; // @[Mux.scala 27:72]
  wire  _T_3092 = btb_rd_addr_f == 8'hc9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1449; // @[Reg.scala 27:20]
  wire [21:0] _T_3403 = _T_3092 ? _T_1449 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3658 = _T_3657 | _T_3403; // @[Mux.scala 27:72]
  wire  _T_3094 = btb_rd_addr_f == 8'hca; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1453; // @[Reg.scala 27:20]
  wire [21:0] _T_3404 = _T_3094 ? _T_1453 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3659 = _T_3658 | _T_3404; // @[Mux.scala 27:72]
  wire  _T_3096 = btb_rd_addr_f == 8'hcb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1457; // @[Reg.scala 27:20]
  wire [21:0] _T_3405 = _T_3096 ? _T_1457 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3660 = _T_3659 | _T_3405; // @[Mux.scala 27:72]
  wire  _T_3098 = btb_rd_addr_f == 8'hcc; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1461; // @[Reg.scala 27:20]
  wire [21:0] _T_3406 = _T_3098 ? _T_1461 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3661 = _T_3660 | _T_3406; // @[Mux.scala 27:72]
  wire  _T_3100 = btb_rd_addr_f == 8'hcd; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1465; // @[Reg.scala 27:20]
  wire [21:0] _T_3407 = _T_3100 ? _T_1465 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3662 = _T_3661 | _T_3407; // @[Mux.scala 27:72]
  wire  _T_3102 = btb_rd_addr_f == 8'hce; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1469; // @[Reg.scala 27:20]
  wire [21:0] _T_3408 = _T_3102 ? _T_1469 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3663 = _T_3662 | _T_3408; // @[Mux.scala 27:72]
  wire  _T_3104 = btb_rd_addr_f == 8'hcf; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1473; // @[Reg.scala 27:20]
  wire [21:0] _T_3409 = _T_3104 ? _T_1473 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3664 = _T_3663 | _T_3409; // @[Mux.scala 27:72]
  wire  _T_3106 = btb_rd_addr_f == 8'hd0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1477; // @[Reg.scala 27:20]
  wire [21:0] _T_3410 = _T_3106 ? _T_1477 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3665 = _T_3664 | _T_3410; // @[Mux.scala 27:72]
  wire  _T_3108 = btb_rd_addr_f == 8'hd1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1481; // @[Reg.scala 27:20]
  wire [21:0] _T_3411 = _T_3108 ? _T_1481 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3666 = _T_3665 | _T_3411; // @[Mux.scala 27:72]
  wire  _T_3110 = btb_rd_addr_f == 8'hd2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1485; // @[Reg.scala 27:20]
  wire [21:0] _T_3412 = _T_3110 ? _T_1485 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3667 = _T_3666 | _T_3412; // @[Mux.scala 27:72]
  wire  _T_3112 = btb_rd_addr_f == 8'hd3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1489; // @[Reg.scala 27:20]
  wire [21:0] _T_3413 = _T_3112 ? _T_1489 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3668 = _T_3667 | _T_3413; // @[Mux.scala 27:72]
  wire  _T_3114 = btb_rd_addr_f == 8'hd4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1493; // @[Reg.scala 27:20]
  wire [21:0] _T_3414 = _T_3114 ? _T_1493 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3669 = _T_3668 | _T_3414; // @[Mux.scala 27:72]
  wire  _T_3116 = btb_rd_addr_f == 8'hd5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1497; // @[Reg.scala 27:20]
  wire [21:0] _T_3415 = _T_3116 ? _T_1497 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3670 = _T_3669 | _T_3415; // @[Mux.scala 27:72]
  wire  _T_3118 = btb_rd_addr_f == 8'hd6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1501; // @[Reg.scala 27:20]
  wire [21:0] _T_3416 = _T_3118 ? _T_1501 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3671 = _T_3670 | _T_3416; // @[Mux.scala 27:72]
  wire  _T_3120 = btb_rd_addr_f == 8'hd7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1505; // @[Reg.scala 27:20]
  wire [21:0] _T_3417 = _T_3120 ? _T_1505 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3672 = _T_3671 | _T_3417; // @[Mux.scala 27:72]
  wire  _T_3122 = btb_rd_addr_f == 8'hd8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1509; // @[Reg.scala 27:20]
  wire [21:0] _T_3418 = _T_3122 ? _T_1509 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3673 = _T_3672 | _T_3418; // @[Mux.scala 27:72]
  wire  _T_3124 = btb_rd_addr_f == 8'hd9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1513; // @[Reg.scala 27:20]
  wire [21:0] _T_3419 = _T_3124 ? _T_1513 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3674 = _T_3673 | _T_3419; // @[Mux.scala 27:72]
  wire  _T_3126 = btb_rd_addr_f == 8'hda; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1517; // @[Reg.scala 27:20]
  wire [21:0] _T_3420 = _T_3126 ? _T_1517 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3675 = _T_3674 | _T_3420; // @[Mux.scala 27:72]
  wire  _T_3128 = btb_rd_addr_f == 8'hdb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1521; // @[Reg.scala 27:20]
  wire [21:0] _T_3421 = _T_3128 ? _T_1521 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3676 = _T_3675 | _T_3421; // @[Mux.scala 27:72]
  wire  _T_3130 = btb_rd_addr_f == 8'hdc; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1525; // @[Reg.scala 27:20]
  wire [21:0] _T_3422 = _T_3130 ? _T_1525 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3677 = _T_3676 | _T_3422; // @[Mux.scala 27:72]
  wire  _T_3132 = btb_rd_addr_f == 8'hdd; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1529; // @[Reg.scala 27:20]
  wire [21:0] _T_3423 = _T_3132 ? _T_1529 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3678 = _T_3677 | _T_3423; // @[Mux.scala 27:72]
  wire  _T_3134 = btb_rd_addr_f == 8'hde; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1533; // @[Reg.scala 27:20]
  wire [21:0] _T_3424 = _T_3134 ? _T_1533 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3679 = _T_3678 | _T_3424; // @[Mux.scala 27:72]
  wire  _T_3136 = btb_rd_addr_f == 8'hdf; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1537; // @[Reg.scala 27:20]
  wire [21:0] _T_3425 = _T_3136 ? _T_1537 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3680 = _T_3679 | _T_3425; // @[Mux.scala 27:72]
  wire  _T_3138 = btb_rd_addr_f == 8'he0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1541; // @[Reg.scala 27:20]
  wire [21:0] _T_3426 = _T_3138 ? _T_1541 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3681 = _T_3680 | _T_3426; // @[Mux.scala 27:72]
  wire  _T_3140 = btb_rd_addr_f == 8'he1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1545; // @[Reg.scala 27:20]
  wire [21:0] _T_3427 = _T_3140 ? _T_1545 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3682 = _T_3681 | _T_3427; // @[Mux.scala 27:72]
  wire  _T_3142 = btb_rd_addr_f == 8'he2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1549; // @[Reg.scala 27:20]
  wire [21:0] _T_3428 = _T_3142 ? _T_1549 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3683 = _T_3682 | _T_3428; // @[Mux.scala 27:72]
  wire  _T_3144 = btb_rd_addr_f == 8'he3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1553; // @[Reg.scala 27:20]
  wire [21:0] _T_3429 = _T_3144 ? _T_1553 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3684 = _T_3683 | _T_3429; // @[Mux.scala 27:72]
  wire  _T_3146 = btb_rd_addr_f == 8'he4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1557; // @[Reg.scala 27:20]
  wire [21:0] _T_3430 = _T_3146 ? _T_1557 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3685 = _T_3684 | _T_3430; // @[Mux.scala 27:72]
  wire  _T_3148 = btb_rd_addr_f == 8'he5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1561; // @[Reg.scala 27:20]
  wire [21:0] _T_3431 = _T_3148 ? _T_1561 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3686 = _T_3685 | _T_3431; // @[Mux.scala 27:72]
  wire  _T_3150 = btb_rd_addr_f == 8'he6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1565; // @[Reg.scala 27:20]
  wire [21:0] _T_3432 = _T_3150 ? _T_1565 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3687 = _T_3686 | _T_3432; // @[Mux.scala 27:72]
  wire  _T_3152 = btb_rd_addr_f == 8'he7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1569; // @[Reg.scala 27:20]
  wire [21:0] _T_3433 = _T_3152 ? _T_1569 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3688 = _T_3687 | _T_3433; // @[Mux.scala 27:72]
  wire  _T_3154 = btb_rd_addr_f == 8'he8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1573; // @[Reg.scala 27:20]
  wire [21:0] _T_3434 = _T_3154 ? _T_1573 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3689 = _T_3688 | _T_3434; // @[Mux.scala 27:72]
  wire  _T_3156 = btb_rd_addr_f == 8'he9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1577; // @[Reg.scala 27:20]
  wire [21:0] _T_3435 = _T_3156 ? _T_1577 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3690 = _T_3689 | _T_3435; // @[Mux.scala 27:72]
  wire  _T_3158 = btb_rd_addr_f == 8'hea; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1581; // @[Reg.scala 27:20]
  wire [21:0] _T_3436 = _T_3158 ? _T_1581 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3691 = _T_3690 | _T_3436; // @[Mux.scala 27:72]
  wire  _T_3160 = btb_rd_addr_f == 8'heb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1585; // @[Reg.scala 27:20]
  wire [21:0] _T_3437 = _T_3160 ? _T_1585 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3692 = _T_3691 | _T_3437; // @[Mux.scala 27:72]
  wire  _T_3162 = btb_rd_addr_f == 8'hec; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1589; // @[Reg.scala 27:20]
  wire [21:0] _T_3438 = _T_3162 ? _T_1589 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3693 = _T_3692 | _T_3438; // @[Mux.scala 27:72]
  wire  _T_3164 = btb_rd_addr_f == 8'hed; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1593; // @[Reg.scala 27:20]
  wire [21:0] _T_3439 = _T_3164 ? _T_1593 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3694 = _T_3693 | _T_3439; // @[Mux.scala 27:72]
  wire  _T_3166 = btb_rd_addr_f == 8'hee; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1597; // @[Reg.scala 27:20]
  wire [21:0] _T_3440 = _T_3166 ? _T_1597 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3695 = _T_3694 | _T_3440; // @[Mux.scala 27:72]
  wire  _T_3168 = btb_rd_addr_f == 8'hef; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1601; // @[Reg.scala 27:20]
  wire [21:0] _T_3441 = _T_3168 ? _T_1601 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3696 = _T_3695 | _T_3441; // @[Mux.scala 27:72]
  wire  _T_3170 = btb_rd_addr_f == 8'hf0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1605; // @[Reg.scala 27:20]
  wire [21:0] _T_3442 = _T_3170 ? _T_1605 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3697 = _T_3696 | _T_3442; // @[Mux.scala 27:72]
  wire  _T_3172 = btb_rd_addr_f == 8'hf1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1609; // @[Reg.scala 27:20]
  wire [21:0] _T_3443 = _T_3172 ? _T_1609 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3698 = _T_3697 | _T_3443; // @[Mux.scala 27:72]
  wire  _T_3174 = btb_rd_addr_f == 8'hf2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1613; // @[Reg.scala 27:20]
  wire [21:0] _T_3444 = _T_3174 ? _T_1613 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3699 = _T_3698 | _T_3444; // @[Mux.scala 27:72]
  wire  _T_3176 = btb_rd_addr_f == 8'hf3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1617; // @[Reg.scala 27:20]
  wire [21:0] _T_3445 = _T_3176 ? _T_1617 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3700 = _T_3699 | _T_3445; // @[Mux.scala 27:72]
  wire  _T_3178 = btb_rd_addr_f == 8'hf4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1621; // @[Reg.scala 27:20]
  wire [21:0] _T_3446 = _T_3178 ? _T_1621 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3701 = _T_3700 | _T_3446; // @[Mux.scala 27:72]
  wire  _T_3180 = btb_rd_addr_f == 8'hf5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1625; // @[Reg.scala 27:20]
  wire [21:0] _T_3447 = _T_3180 ? _T_1625 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3702 = _T_3701 | _T_3447; // @[Mux.scala 27:72]
  wire  _T_3182 = btb_rd_addr_f == 8'hf6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1629; // @[Reg.scala 27:20]
  wire [21:0] _T_3448 = _T_3182 ? _T_1629 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3703 = _T_3702 | _T_3448; // @[Mux.scala 27:72]
  wire  _T_3184 = btb_rd_addr_f == 8'hf7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1633; // @[Reg.scala 27:20]
  wire [21:0] _T_3449 = _T_3184 ? _T_1633 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3704 = _T_3703 | _T_3449; // @[Mux.scala 27:72]
  wire  _T_3186 = btb_rd_addr_f == 8'hf8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1637; // @[Reg.scala 27:20]
  wire [21:0] _T_3450 = _T_3186 ? _T_1637 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3705 = _T_3704 | _T_3450; // @[Mux.scala 27:72]
  wire  _T_3188 = btb_rd_addr_f == 8'hf9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1641; // @[Reg.scala 27:20]
  wire [21:0] _T_3451 = _T_3188 ? _T_1641 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3706 = _T_3705 | _T_3451; // @[Mux.scala 27:72]
  wire  _T_3190 = btb_rd_addr_f == 8'hfa; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1645; // @[Reg.scala 27:20]
  wire [21:0] _T_3452 = _T_3190 ? _T_1645 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3707 = _T_3706 | _T_3452; // @[Mux.scala 27:72]
  wire  _T_3192 = btb_rd_addr_f == 8'hfb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1649; // @[Reg.scala 27:20]
  wire [21:0] _T_3453 = _T_3192 ? _T_1649 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3708 = _T_3707 | _T_3453; // @[Mux.scala 27:72]
  wire  _T_3194 = btb_rd_addr_f == 8'hfc; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1653; // @[Reg.scala 27:20]
  wire [21:0] _T_3454 = _T_3194 ? _T_1653 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3709 = _T_3708 | _T_3454; // @[Mux.scala 27:72]
  wire  _T_3196 = btb_rd_addr_f == 8'hfd; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1657; // @[Reg.scala 27:20]
  wire [21:0] _T_3455 = _T_3196 ? _T_1657 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3710 = _T_3709 | _T_3455; // @[Mux.scala 27:72]
  wire  _T_3198 = btb_rd_addr_f == 8'hfe; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1661; // @[Reg.scala 27:20]
  wire [21:0] _T_3456 = _T_3198 ? _T_1661 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3711 = _T_3710 | _T_3456; // @[Mux.scala 27:72]
  wire  _T_3200 = btb_rd_addr_f == 8'hff; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] _T_1665; // @[Reg.scala 27:20]
  wire [21:0] _T_3457 = _T_3200 ? _T_1665 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3712 = _T_3711 | _T_3457; // @[Mux.scala 27:72]
  wire [21:0] _T_3713 = _T_3712; // @[Mux.scala 27:72 Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_f = _T_3712; // @[ifu_bp_ctl.scala 435:28]
  wire [4:0] _T_29 = io_ifc_fetch_addr_f[13:9] ^ io_ifc_fetch_addr_f[18:14]; // @[lib.scala 42:111]
  wire [4:0] _T_30 = _T_29 ^ io_ifc_fetch_addr_f[23:19]; // @[lib.scala 42:111]
  wire  _T_50 = _T_3713[21:17] == _T_30; // @[ifu_bp_ctl.scala 144:98]
  wire  _T_51 = _T_3713[0] & _T_50; // @[ifu_bp_ctl.scala 144:55]
  wire  _T_19 = io_exu_bp_exu_i0_br_index_r == btb_rd_addr_f; // @[ifu_bp_ctl.scala 125:72]
  wire  branch_error_collision_f = dec_tlu_error_wb & _T_19; // @[ifu_bp_ctl.scala 125:51]
  wire  branch_error_bank_conflict_f = branch_error_collision_f & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 129:63]
  wire  _T_52 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & branch_error_bank_conflict_f; // @[ifu_bp_ctl.scala 145:22]
  wire  _T_53 = ~_T_52; // @[ifu_bp_ctl.scala 145:5]
  wire  _T_54 = _T_51 & _T_53; // @[ifu_bp_ctl.scala 144:118]
  wire  _T_55 = _T_54 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 145:54]
  wire  _T_57 = _T_55 & _T; // @[ifu_bp_ctl.scala 145:75]
  wire  _T_90 = _T_3713[3] ^ _T_3713[4]; // @[ifu_bp_ctl.scala 159:90]
  wire  _T_91 = _T_57 & _T_90; // @[ifu_bp_ctl.scala 159:56]
  wire  _T_95 = ~_T_90; // @[ifu_bp_ctl.scala 160:24]
  wire  _T_96 = _T_57 & _T_95; // @[ifu_bp_ctl.scala 160:22]
  wire [1:0] _T_97 = {_T_91,_T_96}; // @[Cat.scala 29:58]
  wire [21:0] _T_142 = _T_97[1] ? _T_3713 : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] _T_1669; // @[Reg.scala 27:20]
  wire [21:0] _T_4226 = _T_2690 ? _T_1669 : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] _T_1673; // @[Reg.scala 27:20]
  wire [21:0] _T_4227 = _T_2692 ? _T_1673 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4482 = _T_4226 | _T_4227; // @[Mux.scala 27:72]
  reg [21:0] _T_1677; // @[Reg.scala 27:20]
  wire [21:0] _T_4228 = _T_2694 ? _T_1677 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4483 = _T_4482 | _T_4228; // @[Mux.scala 27:72]
  reg [21:0] _T_1681; // @[Reg.scala 27:20]
  wire [21:0] _T_4229 = _T_2696 ? _T_1681 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4484 = _T_4483 | _T_4229; // @[Mux.scala 27:72]
  reg [21:0] _T_1685; // @[Reg.scala 27:20]
  wire [21:0] _T_4230 = _T_2698 ? _T_1685 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4485 = _T_4484 | _T_4230; // @[Mux.scala 27:72]
  reg [21:0] _T_1689; // @[Reg.scala 27:20]
  wire [21:0] _T_4231 = _T_2700 ? _T_1689 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4486 = _T_4485 | _T_4231; // @[Mux.scala 27:72]
  reg [21:0] _T_1693; // @[Reg.scala 27:20]
  wire [21:0] _T_4232 = _T_2702 ? _T_1693 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4487 = _T_4486 | _T_4232; // @[Mux.scala 27:72]
  reg [21:0] _T_1697; // @[Reg.scala 27:20]
  wire [21:0] _T_4233 = _T_2704 ? _T_1697 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4488 = _T_4487 | _T_4233; // @[Mux.scala 27:72]
  reg [21:0] _T_1701; // @[Reg.scala 27:20]
  wire [21:0] _T_4234 = _T_2706 ? _T_1701 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4489 = _T_4488 | _T_4234; // @[Mux.scala 27:72]
  reg [21:0] _T_1705; // @[Reg.scala 27:20]
  wire [21:0] _T_4235 = _T_2708 ? _T_1705 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4490 = _T_4489 | _T_4235; // @[Mux.scala 27:72]
  reg [21:0] _T_1709; // @[Reg.scala 27:20]
  wire [21:0] _T_4236 = _T_2710 ? _T_1709 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4491 = _T_4490 | _T_4236; // @[Mux.scala 27:72]
  reg [21:0] _T_1713; // @[Reg.scala 27:20]
  wire [21:0] _T_4237 = _T_2712 ? _T_1713 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4492 = _T_4491 | _T_4237; // @[Mux.scala 27:72]
  reg [21:0] _T_1717; // @[Reg.scala 27:20]
  wire [21:0] _T_4238 = _T_2714 ? _T_1717 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4493 = _T_4492 | _T_4238; // @[Mux.scala 27:72]
  reg [21:0] _T_1721; // @[Reg.scala 27:20]
  wire [21:0] _T_4239 = _T_2716 ? _T_1721 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4494 = _T_4493 | _T_4239; // @[Mux.scala 27:72]
  reg [21:0] _T_1725; // @[Reg.scala 27:20]
  wire [21:0] _T_4240 = _T_2718 ? _T_1725 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4495 = _T_4494 | _T_4240; // @[Mux.scala 27:72]
  reg [21:0] _T_1729; // @[Reg.scala 27:20]
  wire [21:0] _T_4241 = _T_2720 ? _T_1729 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4496 = _T_4495 | _T_4241; // @[Mux.scala 27:72]
  reg [21:0] _T_1733; // @[Reg.scala 27:20]
  wire [21:0] _T_4242 = _T_2722 ? _T_1733 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4497 = _T_4496 | _T_4242; // @[Mux.scala 27:72]
  reg [21:0] _T_1737; // @[Reg.scala 27:20]
  wire [21:0] _T_4243 = _T_2724 ? _T_1737 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4498 = _T_4497 | _T_4243; // @[Mux.scala 27:72]
  reg [21:0] _T_1741; // @[Reg.scala 27:20]
  wire [21:0] _T_4244 = _T_2726 ? _T_1741 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4499 = _T_4498 | _T_4244; // @[Mux.scala 27:72]
  reg [21:0] _T_1745; // @[Reg.scala 27:20]
  wire [21:0] _T_4245 = _T_2728 ? _T_1745 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4500 = _T_4499 | _T_4245; // @[Mux.scala 27:72]
  reg [21:0] _T_1749; // @[Reg.scala 27:20]
  wire [21:0] _T_4246 = _T_2730 ? _T_1749 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4501 = _T_4500 | _T_4246; // @[Mux.scala 27:72]
  reg [21:0] _T_1753; // @[Reg.scala 27:20]
  wire [21:0] _T_4247 = _T_2732 ? _T_1753 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4502 = _T_4501 | _T_4247; // @[Mux.scala 27:72]
  reg [21:0] _T_1757; // @[Reg.scala 27:20]
  wire [21:0] _T_4248 = _T_2734 ? _T_1757 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4503 = _T_4502 | _T_4248; // @[Mux.scala 27:72]
  reg [21:0] _T_1761; // @[Reg.scala 27:20]
  wire [21:0] _T_4249 = _T_2736 ? _T_1761 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4504 = _T_4503 | _T_4249; // @[Mux.scala 27:72]
  reg [21:0] _T_1765; // @[Reg.scala 27:20]
  wire [21:0] _T_4250 = _T_2738 ? _T_1765 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4505 = _T_4504 | _T_4250; // @[Mux.scala 27:72]
  reg [21:0] _T_1769; // @[Reg.scala 27:20]
  wire [21:0] _T_4251 = _T_2740 ? _T_1769 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4506 = _T_4505 | _T_4251; // @[Mux.scala 27:72]
  reg [21:0] _T_1773; // @[Reg.scala 27:20]
  wire [21:0] _T_4252 = _T_2742 ? _T_1773 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4507 = _T_4506 | _T_4252; // @[Mux.scala 27:72]
  reg [21:0] _T_1777; // @[Reg.scala 27:20]
  wire [21:0] _T_4253 = _T_2744 ? _T_1777 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4508 = _T_4507 | _T_4253; // @[Mux.scala 27:72]
  reg [21:0] _T_1781; // @[Reg.scala 27:20]
  wire [21:0] _T_4254 = _T_2746 ? _T_1781 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4509 = _T_4508 | _T_4254; // @[Mux.scala 27:72]
  reg [21:0] _T_1785; // @[Reg.scala 27:20]
  wire [21:0] _T_4255 = _T_2748 ? _T_1785 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4510 = _T_4509 | _T_4255; // @[Mux.scala 27:72]
  reg [21:0] _T_1789; // @[Reg.scala 27:20]
  wire [21:0] _T_4256 = _T_2750 ? _T_1789 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4511 = _T_4510 | _T_4256; // @[Mux.scala 27:72]
  reg [21:0] _T_1793; // @[Reg.scala 27:20]
  wire [21:0] _T_4257 = _T_2752 ? _T_1793 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4512 = _T_4511 | _T_4257; // @[Mux.scala 27:72]
  reg [21:0] _T_1797; // @[Reg.scala 27:20]
  wire [21:0] _T_4258 = _T_2754 ? _T_1797 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4513 = _T_4512 | _T_4258; // @[Mux.scala 27:72]
  reg [21:0] _T_1801; // @[Reg.scala 27:20]
  wire [21:0] _T_4259 = _T_2756 ? _T_1801 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4514 = _T_4513 | _T_4259; // @[Mux.scala 27:72]
  reg [21:0] _T_1805; // @[Reg.scala 27:20]
  wire [21:0] _T_4260 = _T_2758 ? _T_1805 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4515 = _T_4514 | _T_4260; // @[Mux.scala 27:72]
  reg [21:0] _T_1809; // @[Reg.scala 27:20]
  wire [21:0] _T_4261 = _T_2760 ? _T_1809 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4516 = _T_4515 | _T_4261; // @[Mux.scala 27:72]
  reg [21:0] _T_1813; // @[Reg.scala 27:20]
  wire [21:0] _T_4262 = _T_2762 ? _T_1813 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4517 = _T_4516 | _T_4262; // @[Mux.scala 27:72]
  reg [21:0] _T_1817; // @[Reg.scala 27:20]
  wire [21:0] _T_4263 = _T_2764 ? _T_1817 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4518 = _T_4517 | _T_4263; // @[Mux.scala 27:72]
  reg [21:0] _T_1821; // @[Reg.scala 27:20]
  wire [21:0] _T_4264 = _T_2766 ? _T_1821 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4519 = _T_4518 | _T_4264; // @[Mux.scala 27:72]
  reg [21:0] _T_1825; // @[Reg.scala 27:20]
  wire [21:0] _T_4265 = _T_2768 ? _T_1825 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4520 = _T_4519 | _T_4265; // @[Mux.scala 27:72]
  reg [21:0] _T_1829; // @[Reg.scala 27:20]
  wire [21:0] _T_4266 = _T_2770 ? _T_1829 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4521 = _T_4520 | _T_4266; // @[Mux.scala 27:72]
  reg [21:0] _T_1833; // @[Reg.scala 27:20]
  wire [21:0] _T_4267 = _T_2772 ? _T_1833 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4522 = _T_4521 | _T_4267; // @[Mux.scala 27:72]
  reg [21:0] _T_1837; // @[Reg.scala 27:20]
  wire [21:0] _T_4268 = _T_2774 ? _T_1837 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4523 = _T_4522 | _T_4268; // @[Mux.scala 27:72]
  reg [21:0] _T_1841; // @[Reg.scala 27:20]
  wire [21:0] _T_4269 = _T_2776 ? _T_1841 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4524 = _T_4523 | _T_4269; // @[Mux.scala 27:72]
  reg [21:0] _T_1845; // @[Reg.scala 27:20]
  wire [21:0] _T_4270 = _T_2778 ? _T_1845 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4525 = _T_4524 | _T_4270; // @[Mux.scala 27:72]
  reg [21:0] _T_1849; // @[Reg.scala 27:20]
  wire [21:0] _T_4271 = _T_2780 ? _T_1849 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4526 = _T_4525 | _T_4271; // @[Mux.scala 27:72]
  reg [21:0] _T_1853; // @[Reg.scala 27:20]
  wire [21:0] _T_4272 = _T_2782 ? _T_1853 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4527 = _T_4526 | _T_4272; // @[Mux.scala 27:72]
  reg [21:0] _T_1857; // @[Reg.scala 27:20]
  wire [21:0] _T_4273 = _T_2784 ? _T_1857 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4528 = _T_4527 | _T_4273; // @[Mux.scala 27:72]
  reg [21:0] _T_1861; // @[Reg.scala 27:20]
  wire [21:0] _T_4274 = _T_2786 ? _T_1861 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4529 = _T_4528 | _T_4274; // @[Mux.scala 27:72]
  reg [21:0] _T_1865; // @[Reg.scala 27:20]
  wire [21:0] _T_4275 = _T_2788 ? _T_1865 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4530 = _T_4529 | _T_4275; // @[Mux.scala 27:72]
  reg [21:0] _T_1869; // @[Reg.scala 27:20]
  wire [21:0] _T_4276 = _T_2790 ? _T_1869 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4531 = _T_4530 | _T_4276; // @[Mux.scala 27:72]
  reg [21:0] _T_1873; // @[Reg.scala 27:20]
  wire [21:0] _T_4277 = _T_2792 ? _T_1873 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4532 = _T_4531 | _T_4277; // @[Mux.scala 27:72]
  reg [21:0] _T_1877; // @[Reg.scala 27:20]
  wire [21:0] _T_4278 = _T_2794 ? _T_1877 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4533 = _T_4532 | _T_4278; // @[Mux.scala 27:72]
  reg [21:0] _T_1881; // @[Reg.scala 27:20]
  wire [21:0] _T_4279 = _T_2796 ? _T_1881 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4534 = _T_4533 | _T_4279; // @[Mux.scala 27:72]
  reg [21:0] _T_1885; // @[Reg.scala 27:20]
  wire [21:0] _T_4280 = _T_2798 ? _T_1885 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4535 = _T_4534 | _T_4280; // @[Mux.scala 27:72]
  reg [21:0] _T_1889; // @[Reg.scala 27:20]
  wire [21:0] _T_4281 = _T_2800 ? _T_1889 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4536 = _T_4535 | _T_4281; // @[Mux.scala 27:72]
  reg [21:0] _T_1893; // @[Reg.scala 27:20]
  wire [21:0] _T_4282 = _T_2802 ? _T_1893 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4537 = _T_4536 | _T_4282; // @[Mux.scala 27:72]
  reg [21:0] _T_1897; // @[Reg.scala 27:20]
  wire [21:0] _T_4283 = _T_2804 ? _T_1897 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4538 = _T_4537 | _T_4283; // @[Mux.scala 27:72]
  reg [21:0] _T_1901; // @[Reg.scala 27:20]
  wire [21:0] _T_4284 = _T_2806 ? _T_1901 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4539 = _T_4538 | _T_4284; // @[Mux.scala 27:72]
  reg [21:0] _T_1905; // @[Reg.scala 27:20]
  wire [21:0] _T_4285 = _T_2808 ? _T_1905 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4540 = _T_4539 | _T_4285; // @[Mux.scala 27:72]
  reg [21:0] _T_1909; // @[Reg.scala 27:20]
  wire [21:0] _T_4286 = _T_2810 ? _T_1909 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4541 = _T_4540 | _T_4286; // @[Mux.scala 27:72]
  reg [21:0] _T_1913; // @[Reg.scala 27:20]
  wire [21:0] _T_4287 = _T_2812 ? _T_1913 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4542 = _T_4541 | _T_4287; // @[Mux.scala 27:72]
  reg [21:0] _T_1917; // @[Reg.scala 27:20]
  wire [21:0] _T_4288 = _T_2814 ? _T_1917 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4543 = _T_4542 | _T_4288; // @[Mux.scala 27:72]
  reg [21:0] _T_1921; // @[Reg.scala 27:20]
  wire [21:0] _T_4289 = _T_2816 ? _T_1921 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4544 = _T_4543 | _T_4289; // @[Mux.scala 27:72]
  reg [21:0] _T_1925; // @[Reg.scala 27:20]
  wire [21:0] _T_4290 = _T_2818 ? _T_1925 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4545 = _T_4544 | _T_4290; // @[Mux.scala 27:72]
  reg [21:0] _T_1929; // @[Reg.scala 27:20]
  wire [21:0] _T_4291 = _T_2820 ? _T_1929 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4546 = _T_4545 | _T_4291; // @[Mux.scala 27:72]
  reg [21:0] _T_1933; // @[Reg.scala 27:20]
  wire [21:0] _T_4292 = _T_2822 ? _T_1933 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4547 = _T_4546 | _T_4292; // @[Mux.scala 27:72]
  reg [21:0] _T_1937; // @[Reg.scala 27:20]
  wire [21:0] _T_4293 = _T_2824 ? _T_1937 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4548 = _T_4547 | _T_4293; // @[Mux.scala 27:72]
  reg [21:0] _T_1941; // @[Reg.scala 27:20]
  wire [21:0] _T_4294 = _T_2826 ? _T_1941 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4549 = _T_4548 | _T_4294; // @[Mux.scala 27:72]
  reg [21:0] _T_1945; // @[Reg.scala 27:20]
  wire [21:0] _T_4295 = _T_2828 ? _T_1945 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4550 = _T_4549 | _T_4295; // @[Mux.scala 27:72]
  reg [21:0] _T_1949; // @[Reg.scala 27:20]
  wire [21:0] _T_4296 = _T_2830 ? _T_1949 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4551 = _T_4550 | _T_4296; // @[Mux.scala 27:72]
  reg [21:0] _T_1953; // @[Reg.scala 27:20]
  wire [21:0] _T_4297 = _T_2832 ? _T_1953 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4552 = _T_4551 | _T_4297; // @[Mux.scala 27:72]
  reg [21:0] _T_1957; // @[Reg.scala 27:20]
  wire [21:0] _T_4298 = _T_2834 ? _T_1957 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4553 = _T_4552 | _T_4298; // @[Mux.scala 27:72]
  reg [21:0] _T_1961; // @[Reg.scala 27:20]
  wire [21:0] _T_4299 = _T_2836 ? _T_1961 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4554 = _T_4553 | _T_4299; // @[Mux.scala 27:72]
  reg [21:0] _T_1965; // @[Reg.scala 27:20]
  wire [21:0] _T_4300 = _T_2838 ? _T_1965 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4555 = _T_4554 | _T_4300; // @[Mux.scala 27:72]
  reg [21:0] _T_1969; // @[Reg.scala 27:20]
  wire [21:0] _T_4301 = _T_2840 ? _T_1969 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4556 = _T_4555 | _T_4301; // @[Mux.scala 27:72]
  reg [21:0] _T_1973; // @[Reg.scala 27:20]
  wire [21:0] _T_4302 = _T_2842 ? _T_1973 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4557 = _T_4556 | _T_4302; // @[Mux.scala 27:72]
  reg [21:0] _T_1977; // @[Reg.scala 27:20]
  wire [21:0] _T_4303 = _T_2844 ? _T_1977 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4558 = _T_4557 | _T_4303; // @[Mux.scala 27:72]
  reg [21:0] _T_1981; // @[Reg.scala 27:20]
  wire [21:0] _T_4304 = _T_2846 ? _T_1981 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4559 = _T_4558 | _T_4304; // @[Mux.scala 27:72]
  reg [21:0] _T_1985; // @[Reg.scala 27:20]
  wire [21:0] _T_4305 = _T_2848 ? _T_1985 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4560 = _T_4559 | _T_4305; // @[Mux.scala 27:72]
  reg [21:0] _T_1989; // @[Reg.scala 27:20]
  wire [21:0] _T_4306 = _T_2850 ? _T_1989 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4561 = _T_4560 | _T_4306; // @[Mux.scala 27:72]
  reg [21:0] _T_1993; // @[Reg.scala 27:20]
  wire [21:0] _T_4307 = _T_2852 ? _T_1993 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4562 = _T_4561 | _T_4307; // @[Mux.scala 27:72]
  reg [21:0] _T_1997; // @[Reg.scala 27:20]
  wire [21:0] _T_4308 = _T_2854 ? _T_1997 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4563 = _T_4562 | _T_4308; // @[Mux.scala 27:72]
  reg [21:0] _T_2001; // @[Reg.scala 27:20]
  wire [21:0] _T_4309 = _T_2856 ? _T_2001 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4564 = _T_4563 | _T_4309; // @[Mux.scala 27:72]
  reg [21:0] _T_2005; // @[Reg.scala 27:20]
  wire [21:0] _T_4310 = _T_2858 ? _T_2005 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4565 = _T_4564 | _T_4310; // @[Mux.scala 27:72]
  reg [21:0] _T_2009; // @[Reg.scala 27:20]
  wire [21:0] _T_4311 = _T_2860 ? _T_2009 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4566 = _T_4565 | _T_4311; // @[Mux.scala 27:72]
  reg [21:0] _T_2013; // @[Reg.scala 27:20]
  wire [21:0] _T_4312 = _T_2862 ? _T_2013 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4567 = _T_4566 | _T_4312; // @[Mux.scala 27:72]
  reg [21:0] _T_2017; // @[Reg.scala 27:20]
  wire [21:0] _T_4313 = _T_2864 ? _T_2017 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4568 = _T_4567 | _T_4313; // @[Mux.scala 27:72]
  reg [21:0] _T_2021; // @[Reg.scala 27:20]
  wire [21:0] _T_4314 = _T_2866 ? _T_2021 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4569 = _T_4568 | _T_4314; // @[Mux.scala 27:72]
  reg [21:0] _T_2025; // @[Reg.scala 27:20]
  wire [21:0] _T_4315 = _T_2868 ? _T_2025 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4570 = _T_4569 | _T_4315; // @[Mux.scala 27:72]
  reg [21:0] _T_2029; // @[Reg.scala 27:20]
  wire [21:0] _T_4316 = _T_2870 ? _T_2029 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4571 = _T_4570 | _T_4316; // @[Mux.scala 27:72]
  reg [21:0] _T_2033; // @[Reg.scala 27:20]
  wire [21:0] _T_4317 = _T_2872 ? _T_2033 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4572 = _T_4571 | _T_4317; // @[Mux.scala 27:72]
  reg [21:0] _T_2037; // @[Reg.scala 27:20]
  wire [21:0] _T_4318 = _T_2874 ? _T_2037 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4573 = _T_4572 | _T_4318; // @[Mux.scala 27:72]
  reg [21:0] _T_2041; // @[Reg.scala 27:20]
  wire [21:0] _T_4319 = _T_2876 ? _T_2041 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4574 = _T_4573 | _T_4319; // @[Mux.scala 27:72]
  reg [21:0] _T_2045; // @[Reg.scala 27:20]
  wire [21:0] _T_4320 = _T_2878 ? _T_2045 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4575 = _T_4574 | _T_4320; // @[Mux.scala 27:72]
  reg [21:0] _T_2049; // @[Reg.scala 27:20]
  wire [21:0] _T_4321 = _T_2880 ? _T_2049 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4576 = _T_4575 | _T_4321; // @[Mux.scala 27:72]
  reg [21:0] _T_2053; // @[Reg.scala 27:20]
  wire [21:0] _T_4322 = _T_2882 ? _T_2053 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4577 = _T_4576 | _T_4322; // @[Mux.scala 27:72]
  reg [21:0] _T_2057; // @[Reg.scala 27:20]
  wire [21:0] _T_4323 = _T_2884 ? _T_2057 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4578 = _T_4577 | _T_4323; // @[Mux.scala 27:72]
  reg [21:0] _T_2061; // @[Reg.scala 27:20]
  wire [21:0] _T_4324 = _T_2886 ? _T_2061 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4579 = _T_4578 | _T_4324; // @[Mux.scala 27:72]
  reg [21:0] _T_2065; // @[Reg.scala 27:20]
  wire [21:0] _T_4325 = _T_2888 ? _T_2065 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4580 = _T_4579 | _T_4325; // @[Mux.scala 27:72]
  reg [21:0] _T_2069; // @[Reg.scala 27:20]
  wire [21:0] _T_4326 = _T_2890 ? _T_2069 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4581 = _T_4580 | _T_4326; // @[Mux.scala 27:72]
  reg [21:0] _T_2073; // @[Reg.scala 27:20]
  wire [21:0] _T_4327 = _T_2892 ? _T_2073 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4582 = _T_4581 | _T_4327; // @[Mux.scala 27:72]
  reg [21:0] _T_2077; // @[Reg.scala 27:20]
  wire [21:0] _T_4328 = _T_2894 ? _T_2077 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4583 = _T_4582 | _T_4328; // @[Mux.scala 27:72]
  reg [21:0] _T_2081; // @[Reg.scala 27:20]
  wire [21:0] _T_4329 = _T_2896 ? _T_2081 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4584 = _T_4583 | _T_4329; // @[Mux.scala 27:72]
  reg [21:0] _T_2085; // @[Reg.scala 27:20]
  wire [21:0] _T_4330 = _T_2898 ? _T_2085 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4585 = _T_4584 | _T_4330; // @[Mux.scala 27:72]
  reg [21:0] _T_2089; // @[Reg.scala 27:20]
  wire [21:0] _T_4331 = _T_2900 ? _T_2089 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4586 = _T_4585 | _T_4331; // @[Mux.scala 27:72]
  reg [21:0] _T_2093; // @[Reg.scala 27:20]
  wire [21:0] _T_4332 = _T_2902 ? _T_2093 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4587 = _T_4586 | _T_4332; // @[Mux.scala 27:72]
  reg [21:0] _T_2097; // @[Reg.scala 27:20]
  wire [21:0] _T_4333 = _T_2904 ? _T_2097 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4588 = _T_4587 | _T_4333; // @[Mux.scala 27:72]
  reg [21:0] _T_2101; // @[Reg.scala 27:20]
  wire [21:0] _T_4334 = _T_2906 ? _T_2101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4589 = _T_4588 | _T_4334; // @[Mux.scala 27:72]
  reg [21:0] _T_2105; // @[Reg.scala 27:20]
  wire [21:0] _T_4335 = _T_2908 ? _T_2105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4590 = _T_4589 | _T_4335; // @[Mux.scala 27:72]
  reg [21:0] _T_2109; // @[Reg.scala 27:20]
  wire [21:0] _T_4336 = _T_2910 ? _T_2109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4591 = _T_4590 | _T_4336; // @[Mux.scala 27:72]
  reg [21:0] _T_2113; // @[Reg.scala 27:20]
  wire [21:0] _T_4337 = _T_2912 ? _T_2113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4592 = _T_4591 | _T_4337; // @[Mux.scala 27:72]
  reg [21:0] _T_2117; // @[Reg.scala 27:20]
  wire [21:0] _T_4338 = _T_2914 ? _T_2117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4593 = _T_4592 | _T_4338; // @[Mux.scala 27:72]
  reg [21:0] _T_2121; // @[Reg.scala 27:20]
  wire [21:0] _T_4339 = _T_2916 ? _T_2121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4594 = _T_4593 | _T_4339; // @[Mux.scala 27:72]
  reg [21:0] _T_2125; // @[Reg.scala 27:20]
  wire [21:0] _T_4340 = _T_2918 ? _T_2125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4595 = _T_4594 | _T_4340; // @[Mux.scala 27:72]
  reg [21:0] _T_2129; // @[Reg.scala 27:20]
  wire [21:0] _T_4341 = _T_2920 ? _T_2129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4596 = _T_4595 | _T_4341; // @[Mux.scala 27:72]
  reg [21:0] _T_2133; // @[Reg.scala 27:20]
  wire [21:0] _T_4342 = _T_2922 ? _T_2133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4597 = _T_4596 | _T_4342; // @[Mux.scala 27:72]
  reg [21:0] _T_2137; // @[Reg.scala 27:20]
  wire [21:0] _T_4343 = _T_2924 ? _T_2137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4598 = _T_4597 | _T_4343; // @[Mux.scala 27:72]
  reg [21:0] _T_2141; // @[Reg.scala 27:20]
  wire [21:0] _T_4344 = _T_2926 ? _T_2141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4599 = _T_4598 | _T_4344; // @[Mux.scala 27:72]
  reg [21:0] _T_2145; // @[Reg.scala 27:20]
  wire [21:0] _T_4345 = _T_2928 ? _T_2145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4600 = _T_4599 | _T_4345; // @[Mux.scala 27:72]
  reg [21:0] _T_2149; // @[Reg.scala 27:20]
  wire [21:0] _T_4346 = _T_2930 ? _T_2149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4601 = _T_4600 | _T_4346; // @[Mux.scala 27:72]
  reg [21:0] _T_2153; // @[Reg.scala 27:20]
  wire [21:0] _T_4347 = _T_2932 ? _T_2153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4602 = _T_4601 | _T_4347; // @[Mux.scala 27:72]
  reg [21:0] _T_2157; // @[Reg.scala 27:20]
  wire [21:0] _T_4348 = _T_2934 ? _T_2157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4603 = _T_4602 | _T_4348; // @[Mux.scala 27:72]
  reg [21:0] _T_2161; // @[Reg.scala 27:20]
  wire [21:0] _T_4349 = _T_2936 ? _T_2161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4604 = _T_4603 | _T_4349; // @[Mux.scala 27:72]
  reg [21:0] _T_2165; // @[Reg.scala 27:20]
  wire [21:0] _T_4350 = _T_2938 ? _T_2165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4605 = _T_4604 | _T_4350; // @[Mux.scala 27:72]
  reg [21:0] _T_2169; // @[Reg.scala 27:20]
  wire [21:0] _T_4351 = _T_2940 ? _T_2169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4606 = _T_4605 | _T_4351; // @[Mux.scala 27:72]
  reg [21:0] _T_2173; // @[Reg.scala 27:20]
  wire [21:0] _T_4352 = _T_2942 ? _T_2173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4607 = _T_4606 | _T_4352; // @[Mux.scala 27:72]
  reg [21:0] _T_2177; // @[Reg.scala 27:20]
  wire [21:0] _T_4353 = _T_2944 ? _T_2177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4608 = _T_4607 | _T_4353; // @[Mux.scala 27:72]
  reg [21:0] _T_2181; // @[Reg.scala 27:20]
  wire [21:0] _T_4354 = _T_2946 ? _T_2181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4609 = _T_4608 | _T_4354; // @[Mux.scala 27:72]
  reg [21:0] _T_2185; // @[Reg.scala 27:20]
  wire [21:0] _T_4355 = _T_2948 ? _T_2185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4610 = _T_4609 | _T_4355; // @[Mux.scala 27:72]
  reg [21:0] _T_2189; // @[Reg.scala 27:20]
  wire [21:0] _T_4356 = _T_2950 ? _T_2189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4611 = _T_4610 | _T_4356; // @[Mux.scala 27:72]
  reg [21:0] _T_2193; // @[Reg.scala 27:20]
  wire [21:0] _T_4357 = _T_2952 ? _T_2193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4612 = _T_4611 | _T_4357; // @[Mux.scala 27:72]
  reg [21:0] _T_2197; // @[Reg.scala 27:20]
  wire [21:0] _T_4358 = _T_2954 ? _T_2197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4613 = _T_4612 | _T_4358; // @[Mux.scala 27:72]
  reg [21:0] _T_2201; // @[Reg.scala 27:20]
  wire [21:0] _T_4359 = _T_2956 ? _T_2201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4614 = _T_4613 | _T_4359; // @[Mux.scala 27:72]
  reg [21:0] _T_2205; // @[Reg.scala 27:20]
  wire [21:0] _T_4360 = _T_2958 ? _T_2205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4615 = _T_4614 | _T_4360; // @[Mux.scala 27:72]
  reg [21:0] _T_2209; // @[Reg.scala 27:20]
  wire [21:0] _T_4361 = _T_2960 ? _T_2209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4616 = _T_4615 | _T_4361; // @[Mux.scala 27:72]
  reg [21:0] _T_2213; // @[Reg.scala 27:20]
  wire [21:0] _T_4362 = _T_2962 ? _T_2213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4617 = _T_4616 | _T_4362; // @[Mux.scala 27:72]
  reg [21:0] _T_2217; // @[Reg.scala 27:20]
  wire [21:0] _T_4363 = _T_2964 ? _T_2217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4618 = _T_4617 | _T_4363; // @[Mux.scala 27:72]
  reg [21:0] _T_2221; // @[Reg.scala 27:20]
  wire [21:0] _T_4364 = _T_2966 ? _T_2221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4619 = _T_4618 | _T_4364; // @[Mux.scala 27:72]
  reg [21:0] _T_2225; // @[Reg.scala 27:20]
  wire [21:0] _T_4365 = _T_2968 ? _T_2225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4620 = _T_4619 | _T_4365; // @[Mux.scala 27:72]
  reg [21:0] _T_2229; // @[Reg.scala 27:20]
  wire [21:0] _T_4366 = _T_2970 ? _T_2229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4621 = _T_4620 | _T_4366; // @[Mux.scala 27:72]
  reg [21:0] _T_2233; // @[Reg.scala 27:20]
  wire [21:0] _T_4367 = _T_2972 ? _T_2233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4622 = _T_4621 | _T_4367; // @[Mux.scala 27:72]
  reg [21:0] _T_2237; // @[Reg.scala 27:20]
  wire [21:0] _T_4368 = _T_2974 ? _T_2237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4623 = _T_4622 | _T_4368; // @[Mux.scala 27:72]
  reg [21:0] _T_2241; // @[Reg.scala 27:20]
  wire [21:0] _T_4369 = _T_2976 ? _T_2241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4624 = _T_4623 | _T_4369; // @[Mux.scala 27:72]
  reg [21:0] _T_2245; // @[Reg.scala 27:20]
  wire [21:0] _T_4370 = _T_2978 ? _T_2245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4625 = _T_4624 | _T_4370; // @[Mux.scala 27:72]
  reg [21:0] _T_2249; // @[Reg.scala 27:20]
  wire [21:0] _T_4371 = _T_2980 ? _T_2249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4626 = _T_4625 | _T_4371; // @[Mux.scala 27:72]
  reg [21:0] _T_2253; // @[Reg.scala 27:20]
  wire [21:0] _T_4372 = _T_2982 ? _T_2253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4627 = _T_4626 | _T_4372; // @[Mux.scala 27:72]
  reg [21:0] _T_2257; // @[Reg.scala 27:20]
  wire [21:0] _T_4373 = _T_2984 ? _T_2257 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4628 = _T_4627 | _T_4373; // @[Mux.scala 27:72]
  reg [21:0] _T_2261; // @[Reg.scala 27:20]
  wire [21:0] _T_4374 = _T_2986 ? _T_2261 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4629 = _T_4628 | _T_4374; // @[Mux.scala 27:72]
  reg [21:0] _T_2265; // @[Reg.scala 27:20]
  wire [21:0] _T_4375 = _T_2988 ? _T_2265 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4630 = _T_4629 | _T_4375; // @[Mux.scala 27:72]
  reg [21:0] _T_2269; // @[Reg.scala 27:20]
  wire [21:0] _T_4376 = _T_2990 ? _T_2269 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4631 = _T_4630 | _T_4376; // @[Mux.scala 27:72]
  reg [21:0] _T_2273; // @[Reg.scala 27:20]
  wire [21:0] _T_4377 = _T_2992 ? _T_2273 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4632 = _T_4631 | _T_4377; // @[Mux.scala 27:72]
  reg [21:0] _T_2277; // @[Reg.scala 27:20]
  wire [21:0] _T_4378 = _T_2994 ? _T_2277 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4633 = _T_4632 | _T_4378; // @[Mux.scala 27:72]
  reg [21:0] _T_2281; // @[Reg.scala 27:20]
  wire [21:0] _T_4379 = _T_2996 ? _T_2281 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4634 = _T_4633 | _T_4379; // @[Mux.scala 27:72]
  reg [21:0] _T_2285; // @[Reg.scala 27:20]
  wire [21:0] _T_4380 = _T_2998 ? _T_2285 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4635 = _T_4634 | _T_4380; // @[Mux.scala 27:72]
  reg [21:0] _T_2289; // @[Reg.scala 27:20]
  wire [21:0] _T_4381 = _T_3000 ? _T_2289 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4636 = _T_4635 | _T_4381; // @[Mux.scala 27:72]
  reg [21:0] _T_2293; // @[Reg.scala 27:20]
  wire [21:0] _T_4382 = _T_3002 ? _T_2293 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4637 = _T_4636 | _T_4382; // @[Mux.scala 27:72]
  reg [21:0] _T_2297; // @[Reg.scala 27:20]
  wire [21:0] _T_4383 = _T_3004 ? _T_2297 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4638 = _T_4637 | _T_4383; // @[Mux.scala 27:72]
  reg [21:0] _T_2301; // @[Reg.scala 27:20]
  wire [21:0] _T_4384 = _T_3006 ? _T_2301 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4639 = _T_4638 | _T_4384; // @[Mux.scala 27:72]
  reg [21:0] _T_2305; // @[Reg.scala 27:20]
  wire [21:0] _T_4385 = _T_3008 ? _T_2305 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4640 = _T_4639 | _T_4385; // @[Mux.scala 27:72]
  reg [21:0] _T_2309; // @[Reg.scala 27:20]
  wire [21:0] _T_4386 = _T_3010 ? _T_2309 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4641 = _T_4640 | _T_4386; // @[Mux.scala 27:72]
  reg [21:0] _T_2313; // @[Reg.scala 27:20]
  wire [21:0] _T_4387 = _T_3012 ? _T_2313 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4642 = _T_4641 | _T_4387; // @[Mux.scala 27:72]
  reg [21:0] _T_2317; // @[Reg.scala 27:20]
  wire [21:0] _T_4388 = _T_3014 ? _T_2317 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4643 = _T_4642 | _T_4388; // @[Mux.scala 27:72]
  reg [21:0] _T_2321; // @[Reg.scala 27:20]
  wire [21:0] _T_4389 = _T_3016 ? _T_2321 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4644 = _T_4643 | _T_4389; // @[Mux.scala 27:72]
  reg [21:0] _T_2325; // @[Reg.scala 27:20]
  wire [21:0] _T_4390 = _T_3018 ? _T_2325 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4645 = _T_4644 | _T_4390; // @[Mux.scala 27:72]
  reg [21:0] _T_2329; // @[Reg.scala 27:20]
  wire [21:0] _T_4391 = _T_3020 ? _T_2329 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4646 = _T_4645 | _T_4391; // @[Mux.scala 27:72]
  reg [21:0] _T_2333; // @[Reg.scala 27:20]
  wire [21:0] _T_4392 = _T_3022 ? _T_2333 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4647 = _T_4646 | _T_4392; // @[Mux.scala 27:72]
  reg [21:0] _T_2337; // @[Reg.scala 27:20]
  wire [21:0] _T_4393 = _T_3024 ? _T_2337 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4648 = _T_4647 | _T_4393; // @[Mux.scala 27:72]
  reg [21:0] _T_2341; // @[Reg.scala 27:20]
  wire [21:0] _T_4394 = _T_3026 ? _T_2341 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4649 = _T_4648 | _T_4394; // @[Mux.scala 27:72]
  reg [21:0] _T_2345; // @[Reg.scala 27:20]
  wire [21:0] _T_4395 = _T_3028 ? _T_2345 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4650 = _T_4649 | _T_4395; // @[Mux.scala 27:72]
  reg [21:0] _T_2349; // @[Reg.scala 27:20]
  wire [21:0] _T_4396 = _T_3030 ? _T_2349 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4651 = _T_4650 | _T_4396; // @[Mux.scala 27:72]
  reg [21:0] _T_2353; // @[Reg.scala 27:20]
  wire [21:0] _T_4397 = _T_3032 ? _T_2353 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4652 = _T_4651 | _T_4397; // @[Mux.scala 27:72]
  reg [21:0] _T_2357; // @[Reg.scala 27:20]
  wire [21:0] _T_4398 = _T_3034 ? _T_2357 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4653 = _T_4652 | _T_4398; // @[Mux.scala 27:72]
  reg [21:0] _T_2361; // @[Reg.scala 27:20]
  wire [21:0] _T_4399 = _T_3036 ? _T_2361 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4654 = _T_4653 | _T_4399; // @[Mux.scala 27:72]
  reg [21:0] _T_2365; // @[Reg.scala 27:20]
  wire [21:0] _T_4400 = _T_3038 ? _T_2365 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4655 = _T_4654 | _T_4400; // @[Mux.scala 27:72]
  reg [21:0] _T_2369; // @[Reg.scala 27:20]
  wire [21:0] _T_4401 = _T_3040 ? _T_2369 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4656 = _T_4655 | _T_4401; // @[Mux.scala 27:72]
  reg [21:0] _T_2373; // @[Reg.scala 27:20]
  wire [21:0] _T_4402 = _T_3042 ? _T_2373 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4657 = _T_4656 | _T_4402; // @[Mux.scala 27:72]
  reg [21:0] _T_2377; // @[Reg.scala 27:20]
  wire [21:0] _T_4403 = _T_3044 ? _T_2377 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4658 = _T_4657 | _T_4403; // @[Mux.scala 27:72]
  reg [21:0] _T_2381; // @[Reg.scala 27:20]
  wire [21:0] _T_4404 = _T_3046 ? _T_2381 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4659 = _T_4658 | _T_4404; // @[Mux.scala 27:72]
  reg [21:0] _T_2385; // @[Reg.scala 27:20]
  wire [21:0] _T_4405 = _T_3048 ? _T_2385 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4660 = _T_4659 | _T_4405; // @[Mux.scala 27:72]
  reg [21:0] _T_2389; // @[Reg.scala 27:20]
  wire [21:0] _T_4406 = _T_3050 ? _T_2389 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4661 = _T_4660 | _T_4406; // @[Mux.scala 27:72]
  reg [21:0] _T_2393; // @[Reg.scala 27:20]
  wire [21:0] _T_4407 = _T_3052 ? _T_2393 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4662 = _T_4661 | _T_4407; // @[Mux.scala 27:72]
  reg [21:0] _T_2397; // @[Reg.scala 27:20]
  wire [21:0] _T_4408 = _T_3054 ? _T_2397 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4663 = _T_4662 | _T_4408; // @[Mux.scala 27:72]
  reg [21:0] _T_2401; // @[Reg.scala 27:20]
  wire [21:0] _T_4409 = _T_3056 ? _T_2401 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4664 = _T_4663 | _T_4409; // @[Mux.scala 27:72]
  reg [21:0] _T_2405; // @[Reg.scala 27:20]
  wire [21:0] _T_4410 = _T_3058 ? _T_2405 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4665 = _T_4664 | _T_4410; // @[Mux.scala 27:72]
  reg [21:0] _T_2409; // @[Reg.scala 27:20]
  wire [21:0] _T_4411 = _T_3060 ? _T_2409 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4666 = _T_4665 | _T_4411; // @[Mux.scala 27:72]
  reg [21:0] _T_2413; // @[Reg.scala 27:20]
  wire [21:0] _T_4412 = _T_3062 ? _T_2413 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4667 = _T_4666 | _T_4412; // @[Mux.scala 27:72]
  reg [21:0] _T_2417; // @[Reg.scala 27:20]
  wire [21:0] _T_4413 = _T_3064 ? _T_2417 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4668 = _T_4667 | _T_4413; // @[Mux.scala 27:72]
  reg [21:0] _T_2421; // @[Reg.scala 27:20]
  wire [21:0] _T_4414 = _T_3066 ? _T_2421 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4669 = _T_4668 | _T_4414; // @[Mux.scala 27:72]
  reg [21:0] _T_2425; // @[Reg.scala 27:20]
  wire [21:0] _T_4415 = _T_3068 ? _T_2425 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4670 = _T_4669 | _T_4415; // @[Mux.scala 27:72]
  reg [21:0] _T_2429; // @[Reg.scala 27:20]
  wire [21:0] _T_4416 = _T_3070 ? _T_2429 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4671 = _T_4670 | _T_4416; // @[Mux.scala 27:72]
  reg [21:0] _T_2433; // @[Reg.scala 27:20]
  wire [21:0] _T_4417 = _T_3072 ? _T_2433 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4672 = _T_4671 | _T_4417; // @[Mux.scala 27:72]
  reg [21:0] _T_2437; // @[Reg.scala 27:20]
  wire [21:0] _T_4418 = _T_3074 ? _T_2437 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4673 = _T_4672 | _T_4418; // @[Mux.scala 27:72]
  reg [21:0] _T_2441; // @[Reg.scala 27:20]
  wire [21:0] _T_4419 = _T_3076 ? _T_2441 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4674 = _T_4673 | _T_4419; // @[Mux.scala 27:72]
  reg [21:0] _T_2445; // @[Reg.scala 27:20]
  wire [21:0] _T_4420 = _T_3078 ? _T_2445 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4675 = _T_4674 | _T_4420; // @[Mux.scala 27:72]
  reg [21:0] _T_2449; // @[Reg.scala 27:20]
  wire [21:0] _T_4421 = _T_3080 ? _T_2449 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4676 = _T_4675 | _T_4421; // @[Mux.scala 27:72]
  reg [21:0] _T_2453; // @[Reg.scala 27:20]
  wire [21:0] _T_4422 = _T_3082 ? _T_2453 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4677 = _T_4676 | _T_4422; // @[Mux.scala 27:72]
  reg [21:0] _T_2457; // @[Reg.scala 27:20]
  wire [21:0] _T_4423 = _T_3084 ? _T_2457 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4678 = _T_4677 | _T_4423; // @[Mux.scala 27:72]
  reg [21:0] _T_2461; // @[Reg.scala 27:20]
  wire [21:0] _T_4424 = _T_3086 ? _T_2461 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4679 = _T_4678 | _T_4424; // @[Mux.scala 27:72]
  reg [21:0] _T_2465; // @[Reg.scala 27:20]
  wire [21:0] _T_4425 = _T_3088 ? _T_2465 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4680 = _T_4679 | _T_4425; // @[Mux.scala 27:72]
  reg [21:0] _T_2469; // @[Reg.scala 27:20]
  wire [21:0] _T_4426 = _T_3090 ? _T_2469 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4681 = _T_4680 | _T_4426; // @[Mux.scala 27:72]
  reg [21:0] _T_2473; // @[Reg.scala 27:20]
  wire [21:0] _T_4427 = _T_3092 ? _T_2473 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4682 = _T_4681 | _T_4427; // @[Mux.scala 27:72]
  reg [21:0] _T_2477; // @[Reg.scala 27:20]
  wire [21:0] _T_4428 = _T_3094 ? _T_2477 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4683 = _T_4682 | _T_4428; // @[Mux.scala 27:72]
  reg [21:0] _T_2481; // @[Reg.scala 27:20]
  wire [21:0] _T_4429 = _T_3096 ? _T_2481 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4684 = _T_4683 | _T_4429; // @[Mux.scala 27:72]
  reg [21:0] _T_2485; // @[Reg.scala 27:20]
  wire [21:0] _T_4430 = _T_3098 ? _T_2485 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4685 = _T_4684 | _T_4430; // @[Mux.scala 27:72]
  reg [21:0] _T_2489; // @[Reg.scala 27:20]
  wire [21:0] _T_4431 = _T_3100 ? _T_2489 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4686 = _T_4685 | _T_4431; // @[Mux.scala 27:72]
  reg [21:0] _T_2493; // @[Reg.scala 27:20]
  wire [21:0] _T_4432 = _T_3102 ? _T_2493 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4687 = _T_4686 | _T_4432; // @[Mux.scala 27:72]
  reg [21:0] _T_2497; // @[Reg.scala 27:20]
  wire [21:0] _T_4433 = _T_3104 ? _T_2497 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4688 = _T_4687 | _T_4433; // @[Mux.scala 27:72]
  reg [21:0] _T_2501; // @[Reg.scala 27:20]
  wire [21:0] _T_4434 = _T_3106 ? _T_2501 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4689 = _T_4688 | _T_4434; // @[Mux.scala 27:72]
  reg [21:0] _T_2505; // @[Reg.scala 27:20]
  wire [21:0] _T_4435 = _T_3108 ? _T_2505 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4690 = _T_4689 | _T_4435; // @[Mux.scala 27:72]
  reg [21:0] _T_2509; // @[Reg.scala 27:20]
  wire [21:0] _T_4436 = _T_3110 ? _T_2509 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4691 = _T_4690 | _T_4436; // @[Mux.scala 27:72]
  reg [21:0] _T_2513; // @[Reg.scala 27:20]
  wire [21:0] _T_4437 = _T_3112 ? _T_2513 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4692 = _T_4691 | _T_4437; // @[Mux.scala 27:72]
  reg [21:0] _T_2517; // @[Reg.scala 27:20]
  wire [21:0] _T_4438 = _T_3114 ? _T_2517 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4693 = _T_4692 | _T_4438; // @[Mux.scala 27:72]
  reg [21:0] _T_2521; // @[Reg.scala 27:20]
  wire [21:0] _T_4439 = _T_3116 ? _T_2521 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4694 = _T_4693 | _T_4439; // @[Mux.scala 27:72]
  reg [21:0] _T_2525; // @[Reg.scala 27:20]
  wire [21:0] _T_4440 = _T_3118 ? _T_2525 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4695 = _T_4694 | _T_4440; // @[Mux.scala 27:72]
  reg [21:0] _T_2529; // @[Reg.scala 27:20]
  wire [21:0] _T_4441 = _T_3120 ? _T_2529 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4696 = _T_4695 | _T_4441; // @[Mux.scala 27:72]
  reg [21:0] _T_2533; // @[Reg.scala 27:20]
  wire [21:0] _T_4442 = _T_3122 ? _T_2533 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4697 = _T_4696 | _T_4442; // @[Mux.scala 27:72]
  reg [21:0] _T_2537; // @[Reg.scala 27:20]
  wire [21:0] _T_4443 = _T_3124 ? _T_2537 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4698 = _T_4697 | _T_4443; // @[Mux.scala 27:72]
  reg [21:0] _T_2541; // @[Reg.scala 27:20]
  wire [21:0] _T_4444 = _T_3126 ? _T_2541 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4699 = _T_4698 | _T_4444; // @[Mux.scala 27:72]
  reg [21:0] _T_2545; // @[Reg.scala 27:20]
  wire [21:0] _T_4445 = _T_3128 ? _T_2545 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4700 = _T_4699 | _T_4445; // @[Mux.scala 27:72]
  reg [21:0] _T_2549; // @[Reg.scala 27:20]
  wire [21:0] _T_4446 = _T_3130 ? _T_2549 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4701 = _T_4700 | _T_4446; // @[Mux.scala 27:72]
  reg [21:0] _T_2553; // @[Reg.scala 27:20]
  wire [21:0] _T_4447 = _T_3132 ? _T_2553 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4702 = _T_4701 | _T_4447; // @[Mux.scala 27:72]
  reg [21:0] _T_2557; // @[Reg.scala 27:20]
  wire [21:0] _T_4448 = _T_3134 ? _T_2557 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4703 = _T_4702 | _T_4448; // @[Mux.scala 27:72]
  reg [21:0] _T_2561; // @[Reg.scala 27:20]
  wire [21:0] _T_4449 = _T_3136 ? _T_2561 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4704 = _T_4703 | _T_4449; // @[Mux.scala 27:72]
  reg [21:0] _T_2565; // @[Reg.scala 27:20]
  wire [21:0] _T_4450 = _T_3138 ? _T_2565 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4705 = _T_4704 | _T_4450; // @[Mux.scala 27:72]
  reg [21:0] _T_2569; // @[Reg.scala 27:20]
  wire [21:0] _T_4451 = _T_3140 ? _T_2569 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4706 = _T_4705 | _T_4451; // @[Mux.scala 27:72]
  reg [21:0] _T_2573; // @[Reg.scala 27:20]
  wire [21:0] _T_4452 = _T_3142 ? _T_2573 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4707 = _T_4706 | _T_4452; // @[Mux.scala 27:72]
  reg [21:0] _T_2577; // @[Reg.scala 27:20]
  wire [21:0] _T_4453 = _T_3144 ? _T_2577 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4708 = _T_4707 | _T_4453; // @[Mux.scala 27:72]
  reg [21:0] _T_2581; // @[Reg.scala 27:20]
  wire [21:0] _T_4454 = _T_3146 ? _T_2581 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4709 = _T_4708 | _T_4454; // @[Mux.scala 27:72]
  reg [21:0] _T_2585; // @[Reg.scala 27:20]
  wire [21:0] _T_4455 = _T_3148 ? _T_2585 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4710 = _T_4709 | _T_4455; // @[Mux.scala 27:72]
  reg [21:0] _T_2589; // @[Reg.scala 27:20]
  wire [21:0] _T_4456 = _T_3150 ? _T_2589 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4711 = _T_4710 | _T_4456; // @[Mux.scala 27:72]
  reg [21:0] _T_2593; // @[Reg.scala 27:20]
  wire [21:0] _T_4457 = _T_3152 ? _T_2593 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4712 = _T_4711 | _T_4457; // @[Mux.scala 27:72]
  reg [21:0] _T_2597; // @[Reg.scala 27:20]
  wire [21:0] _T_4458 = _T_3154 ? _T_2597 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4713 = _T_4712 | _T_4458; // @[Mux.scala 27:72]
  reg [21:0] _T_2601; // @[Reg.scala 27:20]
  wire [21:0] _T_4459 = _T_3156 ? _T_2601 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4714 = _T_4713 | _T_4459; // @[Mux.scala 27:72]
  reg [21:0] _T_2605; // @[Reg.scala 27:20]
  wire [21:0] _T_4460 = _T_3158 ? _T_2605 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4715 = _T_4714 | _T_4460; // @[Mux.scala 27:72]
  reg [21:0] _T_2609; // @[Reg.scala 27:20]
  wire [21:0] _T_4461 = _T_3160 ? _T_2609 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4716 = _T_4715 | _T_4461; // @[Mux.scala 27:72]
  reg [21:0] _T_2613; // @[Reg.scala 27:20]
  wire [21:0] _T_4462 = _T_3162 ? _T_2613 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4717 = _T_4716 | _T_4462; // @[Mux.scala 27:72]
  reg [21:0] _T_2617; // @[Reg.scala 27:20]
  wire [21:0] _T_4463 = _T_3164 ? _T_2617 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4718 = _T_4717 | _T_4463; // @[Mux.scala 27:72]
  reg [21:0] _T_2621; // @[Reg.scala 27:20]
  wire [21:0] _T_4464 = _T_3166 ? _T_2621 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4719 = _T_4718 | _T_4464; // @[Mux.scala 27:72]
  reg [21:0] _T_2625; // @[Reg.scala 27:20]
  wire [21:0] _T_4465 = _T_3168 ? _T_2625 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4720 = _T_4719 | _T_4465; // @[Mux.scala 27:72]
  reg [21:0] _T_2629; // @[Reg.scala 27:20]
  wire [21:0] _T_4466 = _T_3170 ? _T_2629 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4721 = _T_4720 | _T_4466; // @[Mux.scala 27:72]
  reg [21:0] _T_2633; // @[Reg.scala 27:20]
  wire [21:0] _T_4467 = _T_3172 ? _T_2633 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4722 = _T_4721 | _T_4467; // @[Mux.scala 27:72]
  reg [21:0] _T_2637; // @[Reg.scala 27:20]
  wire [21:0] _T_4468 = _T_3174 ? _T_2637 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4723 = _T_4722 | _T_4468; // @[Mux.scala 27:72]
  reg [21:0] _T_2641; // @[Reg.scala 27:20]
  wire [21:0] _T_4469 = _T_3176 ? _T_2641 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4724 = _T_4723 | _T_4469; // @[Mux.scala 27:72]
  reg [21:0] _T_2645; // @[Reg.scala 27:20]
  wire [21:0] _T_4470 = _T_3178 ? _T_2645 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4725 = _T_4724 | _T_4470; // @[Mux.scala 27:72]
  reg [21:0] _T_2649; // @[Reg.scala 27:20]
  wire [21:0] _T_4471 = _T_3180 ? _T_2649 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4726 = _T_4725 | _T_4471; // @[Mux.scala 27:72]
  reg [21:0] _T_2653; // @[Reg.scala 27:20]
  wire [21:0] _T_4472 = _T_3182 ? _T_2653 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4727 = _T_4726 | _T_4472; // @[Mux.scala 27:72]
  reg [21:0] _T_2657; // @[Reg.scala 27:20]
  wire [21:0] _T_4473 = _T_3184 ? _T_2657 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4728 = _T_4727 | _T_4473; // @[Mux.scala 27:72]
  reg [21:0] _T_2661; // @[Reg.scala 27:20]
  wire [21:0] _T_4474 = _T_3186 ? _T_2661 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4729 = _T_4728 | _T_4474; // @[Mux.scala 27:72]
  reg [21:0] _T_2665; // @[Reg.scala 27:20]
  wire [21:0] _T_4475 = _T_3188 ? _T_2665 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4730 = _T_4729 | _T_4475; // @[Mux.scala 27:72]
  reg [21:0] _T_2669; // @[Reg.scala 27:20]
  wire [21:0] _T_4476 = _T_3190 ? _T_2669 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4731 = _T_4730 | _T_4476; // @[Mux.scala 27:72]
  reg [21:0] _T_2673; // @[Reg.scala 27:20]
  wire [21:0] _T_4477 = _T_3192 ? _T_2673 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4732 = _T_4731 | _T_4477; // @[Mux.scala 27:72]
  reg [21:0] _T_2677; // @[Reg.scala 27:20]
  wire [21:0] _T_4478 = _T_3194 ? _T_2677 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4733 = _T_4732 | _T_4478; // @[Mux.scala 27:72]
  reg [21:0] _T_2681; // @[Reg.scala 27:20]
  wire [21:0] _T_4479 = _T_3196 ? _T_2681 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4734 = _T_4733 | _T_4479; // @[Mux.scala 27:72]
  reg [21:0] _T_2685; // @[Reg.scala 27:20]
  wire [21:0] _T_4480 = _T_3198 ? _T_2685 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4735 = _T_4734 | _T_4480; // @[Mux.scala 27:72]
  reg [21:0] _T_2689; // @[Reg.scala 27:20]
  wire [21:0] _T_4481 = _T_3200 ? _T_2689 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4736 = _T_4735 | _T_4481; // @[Mux.scala 27:72]
  wire [21:0] _T_4737 = _T_4736; // @[Mux.scala 27:72 Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_f = _T_4736; // @[ifu_bp_ctl.scala 438:28]
  wire  _T_60 = _T_4737[21:17] == _T_30; // @[ifu_bp_ctl.scala 148:98]
  wire  _T_61 = _T_4737[0] & _T_60; // @[ifu_bp_ctl.scala 148:55]
  wire  _T_64 = _T_61 & _T_53; // @[ifu_bp_ctl.scala 148:118]
  wire  _T_65 = _T_64 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 149:54]
  wire  _T_67 = _T_65 & _T; // @[ifu_bp_ctl.scala 149:75]
  wire  _T_100 = _T_4737[3] ^ _T_4737[4]; // @[ifu_bp_ctl.scala 162:90]
  wire  _T_101 = _T_67 & _T_100; // @[ifu_bp_ctl.scala 162:56]
  wire  _T_105 = ~_T_100; // @[ifu_bp_ctl.scala 163:24]
  wire  _T_106 = _T_67 & _T_105; // @[ifu_bp_ctl.scala 163:22]
  wire [1:0] _T_107 = {_T_101,_T_106}; // @[Cat.scala 29:58]
  wire [21:0] _T_143 = _T_107[1] ? _T_4737 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_144 = _T_142 | _T_143; // @[Mux.scala 27:72]
  wire [21:0] _T_164 = _T_162 ? _T_144 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4738 = btb_rd_addr_p1_f == 8'h0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5250 = _T_4738 ? _T_645 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4740 = btb_rd_addr_p1_f == 8'h1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5251 = _T_4740 ? _T_649 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5506 = _T_5250 | _T_5251; // @[Mux.scala 27:72]
  wire  _T_4742 = btb_rd_addr_p1_f == 8'h2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5252 = _T_4742 ? _T_653 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5507 = _T_5506 | _T_5252; // @[Mux.scala 27:72]
  wire  _T_4744 = btb_rd_addr_p1_f == 8'h3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5253 = _T_4744 ? _T_657 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5508 = _T_5507 | _T_5253; // @[Mux.scala 27:72]
  wire  _T_4746 = btb_rd_addr_p1_f == 8'h4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5254 = _T_4746 ? _T_661 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5509 = _T_5508 | _T_5254; // @[Mux.scala 27:72]
  wire  _T_4748 = btb_rd_addr_p1_f == 8'h5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5255 = _T_4748 ? _T_665 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5510 = _T_5509 | _T_5255; // @[Mux.scala 27:72]
  wire  _T_4750 = btb_rd_addr_p1_f == 8'h6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5256 = _T_4750 ? _T_669 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5511 = _T_5510 | _T_5256; // @[Mux.scala 27:72]
  wire  _T_4752 = btb_rd_addr_p1_f == 8'h7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5257 = _T_4752 ? _T_673 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5512 = _T_5511 | _T_5257; // @[Mux.scala 27:72]
  wire  _T_4754 = btb_rd_addr_p1_f == 8'h8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5258 = _T_4754 ? _T_677 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5513 = _T_5512 | _T_5258; // @[Mux.scala 27:72]
  wire  _T_4756 = btb_rd_addr_p1_f == 8'h9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5259 = _T_4756 ? _T_681 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5514 = _T_5513 | _T_5259; // @[Mux.scala 27:72]
  wire  _T_4758 = btb_rd_addr_p1_f == 8'ha; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5260 = _T_4758 ? _T_685 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5515 = _T_5514 | _T_5260; // @[Mux.scala 27:72]
  wire  _T_4760 = btb_rd_addr_p1_f == 8'hb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5261 = _T_4760 ? _T_689 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5516 = _T_5515 | _T_5261; // @[Mux.scala 27:72]
  wire  _T_4762 = btb_rd_addr_p1_f == 8'hc; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5262 = _T_4762 ? _T_693 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5517 = _T_5516 | _T_5262; // @[Mux.scala 27:72]
  wire  _T_4764 = btb_rd_addr_p1_f == 8'hd; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5263 = _T_4764 ? _T_697 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5518 = _T_5517 | _T_5263; // @[Mux.scala 27:72]
  wire  _T_4766 = btb_rd_addr_p1_f == 8'he; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5264 = _T_4766 ? _T_701 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5519 = _T_5518 | _T_5264; // @[Mux.scala 27:72]
  wire  _T_4768 = btb_rd_addr_p1_f == 8'hf; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5265 = _T_4768 ? _T_705 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5520 = _T_5519 | _T_5265; // @[Mux.scala 27:72]
  wire  _T_4770 = btb_rd_addr_p1_f == 8'h10; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5266 = _T_4770 ? _T_709 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5521 = _T_5520 | _T_5266; // @[Mux.scala 27:72]
  wire  _T_4772 = btb_rd_addr_p1_f == 8'h11; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5267 = _T_4772 ? _T_713 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5522 = _T_5521 | _T_5267; // @[Mux.scala 27:72]
  wire  _T_4774 = btb_rd_addr_p1_f == 8'h12; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5268 = _T_4774 ? _T_717 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5523 = _T_5522 | _T_5268; // @[Mux.scala 27:72]
  wire  _T_4776 = btb_rd_addr_p1_f == 8'h13; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5269 = _T_4776 ? _T_721 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5524 = _T_5523 | _T_5269; // @[Mux.scala 27:72]
  wire  _T_4778 = btb_rd_addr_p1_f == 8'h14; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5270 = _T_4778 ? _T_725 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5525 = _T_5524 | _T_5270; // @[Mux.scala 27:72]
  wire  _T_4780 = btb_rd_addr_p1_f == 8'h15; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5271 = _T_4780 ? _T_729 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5526 = _T_5525 | _T_5271; // @[Mux.scala 27:72]
  wire  _T_4782 = btb_rd_addr_p1_f == 8'h16; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5272 = _T_4782 ? _T_733 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5527 = _T_5526 | _T_5272; // @[Mux.scala 27:72]
  wire  _T_4784 = btb_rd_addr_p1_f == 8'h17; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5273 = _T_4784 ? _T_737 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5528 = _T_5527 | _T_5273; // @[Mux.scala 27:72]
  wire  _T_4786 = btb_rd_addr_p1_f == 8'h18; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5274 = _T_4786 ? _T_741 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5529 = _T_5528 | _T_5274; // @[Mux.scala 27:72]
  wire  _T_4788 = btb_rd_addr_p1_f == 8'h19; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5275 = _T_4788 ? _T_745 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5530 = _T_5529 | _T_5275; // @[Mux.scala 27:72]
  wire  _T_4790 = btb_rd_addr_p1_f == 8'h1a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5276 = _T_4790 ? _T_749 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5531 = _T_5530 | _T_5276; // @[Mux.scala 27:72]
  wire  _T_4792 = btb_rd_addr_p1_f == 8'h1b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5277 = _T_4792 ? _T_753 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5532 = _T_5531 | _T_5277; // @[Mux.scala 27:72]
  wire  _T_4794 = btb_rd_addr_p1_f == 8'h1c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5278 = _T_4794 ? _T_757 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5533 = _T_5532 | _T_5278; // @[Mux.scala 27:72]
  wire  _T_4796 = btb_rd_addr_p1_f == 8'h1d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5279 = _T_4796 ? _T_761 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5534 = _T_5533 | _T_5279; // @[Mux.scala 27:72]
  wire  _T_4798 = btb_rd_addr_p1_f == 8'h1e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5280 = _T_4798 ? _T_765 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5535 = _T_5534 | _T_5280; // @[Mux.scala 27:72]
  wire  _T_4800 = btb_rd_addr_p1_f == 8'h1f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5281 = _T_4800 ? _T_769 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5536 = _T_5535 | _T_5281; // @[Mux.scala 27:72]
  wire  _T_4802 = btb_rd_addr_p1_f == 8'h20; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5282 = _T_4802 ? _T_773 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5537 = _T_5536 | _T_5282; // @[Mux.scala 27:72]
  wire  _T_4804 = btb_rd_addr_p1_f == 8'h21; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5283 = _T_4804 ? _T_777 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5538 = _T_5537 | _T_5283; // @[Mux.scala 27:72]
  wire  _T_4806 = btb_rd_addr_p1_f == 8'h22; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5284 = _T_4806 ? _T_781 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5539 = _T_5538 | _T_5284; // @[Mux.scala 27:72]
  wire  _T_4808 = btb_rd_addr_p1_f == 8'h23; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5285 = _T_4808 ? _T_785 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5540 = _T_5539 | _T_5285; // @[Mux.scala 27:72]
  wire  _T_4810 = btb_rd_addr_p1_f == 8'h24; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5286 = _T_4810 ? _T_789 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5541 = _T_5540 | _T_5286; // @[Mux.scala 27:72]
  wire  _T_4812 = btb_rd_addr_p1_f == 8'h25; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5287 = _T_4812 ? _T_793 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5542 = _T_5541 | _T_5287; // @[Mux.scala 27:72]
  wire  _T_4814 = btb_rd_addr_p1_f == 8'h26; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5288 = _T_4814 ? _T_797 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5543 = _T_5542 | _T_5288; // @[Mux.scala 27:72]
  wire  _T_4816 = btb_rd_addr_p1_f == 8'h27; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5289 = _T_4816 ? _T_801 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5544 = _T_5543 | _T_5289; // @[Mux.scala 27:72]
  wire  _T_4818 = btb_rd_addr_p1_f == 8'h28; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5290 = _T_4818 ? _T_805 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5545 = _T_5544 | _T_5290; // @[Mux.scala 27:72]
  wire  _T_4820 = btb_rd_addr_p1_f == 8'h29; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5291 = _T_4820 ? _T_809 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5546 = _T_5545 | _T_5291; // @[Mux.scala 27:72]
  wire  _T_4822 = btb_rd_addr_p1_f == 8'h2a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5292 = _T_4822 ? _T_813 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5547 = _T_5546 | _T_5292; // @[Mux.scala 27:72]
  wire  _T_4824 = btb_rd_addr_p1_f == 8'h2b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5293 = _T_4824 ? _T_817 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5548 = _T_5547 | _T_5293; // @[Mux.scala 27:72]
  wire  _T_4826 = btb_rd_addr_p1_f == 8'h2c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5294 = _T_4826 ? _T_821 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5549 = _T_5548 | _T_5294; // @[Mux.scala 27:72]
  wire  _T_4828 = btb_rd_addr_p1_f == 8'h2d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5295 = _T_4828 ? _T_825 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5550 = _T_5549 | _T_5295; // @[Mux.scala 27:72]
  wire  _T_4830 = btb_rd_addr_p1_f == 8'h2e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5296 = _T_4830 ? _T_829 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5551 = _T_5550 | _T_5296; // @[Mux.scala 27:72]
  wire  _T_4832 = btb_rd_addr_p1_f == 8'h2f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5297 = _T_4832 ? _T_833 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5552 = _T_5551 | _T_5297; // @[Mux.scala 27:72]
  wire  _T_4834 = btb_rd_addr_p1_f == 8'h30; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5298 = _T_4834 ? _T_837 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5553 = _T_5552 | _T_5298; // @[Mux.scala 27:72]
  wire  _T_4836 = btb_rd_addr_p1_f == 8'h31; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5299 = _T_4836 ? _T_841 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5554 = _T_5553 | _T_5299; // @[Mux.scala 27:72]
  wire  _T_4838 = btb_rd_addr_p1_f == 8'h32; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5300 = _T_4838 ? _T_845 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5555 = _T_5554 | _T_5300; // @[Mux.scala 27:72]
  wire  _T_4840 = btb_rd_addr_p1_f == 8'h33; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5301 = _T_4840 ? _T_849 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5556 = _T_5555 | _T_5301; // @[Mux.scala 27:72]
  wire  _T_4842 = btb_rd_addr_p1_f == 8'h34; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5302 = _T_4842 ? _T_853 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5557 = _T_5556 | _T_5302; // @[Mux.scala 27:72]
  wire  _T_4844 = btb_rd_addr_p1_f == 8'h35; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5303 = _T_4844 ? _T_857 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5558 = _T_5557 | _T_5303; // @[Mux.scala 27:72]
  wire  _T_4846 = btb_rd_addr_p1_f == 8'h36; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5304 = _T_4846 ? _T_861 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5559 = _T_5558 | _T_5304; // @[Mux.scala 27:72]
  wire  _T_4848 = btb_rd_addr_p1_f == 8'h37; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5305 = _T_4848 ? _T_865 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5560 = _T_5559 | _T_5305; // @[Mux.scala 27:72]
  wire  _T_4850 = btb_rd_addr_p1_f == 8'h38; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5306 = _T_4850 ? _T_869 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5561 = _T_5560 | _T_5306; // @[Mux.scala 27:72]
  wire  _T_4852 = btb_rd_addr_p1_f == 8'h39; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5307 = _T_4852 ? _T_873 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5562 = _T_5561 | _T_5307; // @[Mux.scala 27:72]
  wire  _T_4854 = btb_rd_addr_p1_f == 8'h3a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5308 = _T_4854 ? _T_877 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5563 = _T_5562 | _T_5308; // @[Mux.scala 27:72]
  wire  _T_4856 = btb_rd_addr_p1_f == 8'h3b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5309 = _T_4856 ? _T_881 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5564 = _T_5563 | _T_5309; // @[Mux.scala 27:72]
  wire  _T_4858 = btb_rd_addr_p1_f == 8'h3c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5310 = _T_4858 ? _T_885 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5565 = _T_5564 | _T_5310; // @[Mux.scala 27:72]
  wire  _T_4860 = btb_rd_addr_p1_f == 8'h3d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5311 = _T_4860 ? _T_889 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5566 = _T_5565 | _T_5311; // @[Mux.scala 27:72]
  wire  _T_4862 = btb_rd_addr_p1_f == 8'h3e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5312 = _T_4862 ? _T_893 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5567 = _T_5566 | _T_5312; // @[Mux.scala 27:72]
  wire  _T_4864 = btb_rd_addr_p1_f == 8'h3f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5313 = _T_4864 ? _T_897 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5568 = _T_5567 | _T_5313; // @[Mux.scala 27:72]
  wire  _T_4866 = btb_rd_addr_p1_f == 8'h40; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5314 = _T_4866 ? _T_901 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5569 = _T_5568 | _T_5314; // @[Mux.scala 27:72]
  wire  _T_4868 = btb_rd_addr_p1_f == 8'h41; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5315 = _T_4868 ? _T_905 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5570 = _T_5569 | _T_5315; // @[Mux.scala 27:72]
  wire  _T_4870 = btb_rd_addr_p1_f == 8'h42; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5316 = _T_4870 ? _T_909 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5571 = _T_5570 | _T_5316; // @[Mux.scala 27:72]
  wire  _T_4872 = btb_rd_addr_p1_f == 8'h43; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5317 = _T_4872 ? _T_913 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5572 = _T_5571 | _T_5317; // @[Mux.scala 27:72]
  wire  _T_4874 = btb_rd_addr_p1_f == 8'h44; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5318 = _T_4874 ? _T_917 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5573 = _T_5572 | _T_5318; // @[Mux.scala 27:72]
  wire  _T_4876 = btb_rd_addr_p1_f == 8'h45; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5319 = _T_4876 ? _T_921 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5574 = _T_5573 | _T_5319; // @[Mux.scala 27:72]
  wire  _T_4878 = btb_rd_addr_p1_f == 8'h46; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5320 = _T_4878 ? _T_925 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5575 = _T_5574 | _T_5320; // @[Mux.scala 27:72]
  wire  _T_4880 = btb_rd_addr_p1_f == 8'h47; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5321 = _T_4880 ? _T_929 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5576 = _T_5575 | _T_5321; // @[Mux.scala 27:72]
  wire  _T_4882 = btb_rd_addr_p1_f == 8'h48; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5322 = _T_4882 ? _T_933 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5577 = _T_5576 | _T_5322; // @[Mux.scala 27:72]
  wire  _T_4884 = btb_rd_addr_p1_f == 8'h49; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5323 = _T_4884 ? _T_937 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5578 = _T_5577 | _T_5323; // @[Mux.scala 27:72]
  wire  _T_4886 = btb_rd_addr_p1_f == 8'h4a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5324 = _T_4886 ? _T_941 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5579 = _T_5578 | _T_5324; // @[Mux.scala 27:72]
  wire  _T_4888 = btb_rd_addr_p1_f == 8'h4b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5325 = _T_4888 ? _T_945 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5580 = _T_5579 | _T_5325; // @[Mux.scala 27:72]
  wire  _T_4890 = btb_rd_addr_p1_f == 8'h4c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5326 = _T_4890 ? _T_949 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5581 = _T_5580 | _T_5326; // @[Mux.scala 27:72]
  wire  _T_4892 = btb_rd_addr_p1_f == 8'h4d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5327 = _T_4892 ? _T_953 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5582 = _T_5581 | _T_5327; // @[Mux.scala 27:72]
  wire  _T_4894 = btb_rd_addr_p1_f == 8'h4e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5328 = _T_4894 ? _T_957 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5583 = _T_5582 | _T_5328; // @[Mux.scala 27:72]
  wire  _T_4896 = btb_rd_addr_p1_f == 8'h4f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5329 = _T_4896 ? _T_961 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5584 = _T_5583 | _T_5329; // @[Mux.scala 27:72]
  wire  _T_4898 = btb_rd_addr_p1_f == 8'h50; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5330 = _T_4898 ? _T_965 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5585 = _T_5584 | _T_5330; // @[Mux.scala 27:72]
  wire  _T_4900 = btb_rd_addr_p1_f == 8'h51; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5331 = _T_4900 ? _T_969 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5586 = _T_5585 | _T_5331; // @[Mux.scala 27:72]
  wire  _T_4902 = btb_rd_addr_p1_f == 8'h52; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5332 = _T_4902 ? _T_973 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5587 = _T_5586 | _T_5332; // @[Mux.scala 27:72]
  wire  _T_4904 = btb_rd_addr_p1_f == 8'h53; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5333 = _T_4904 ? _T_977 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5588 = _T_5587 | _T_5333; // @[Mux.scala 27:72]
  wire  _T_4906 = btb_rd_addr_p1_f == 8'h54; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5334 = _T_4906 ? _T_981 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5589 = _T_5588 | _T_5334; // @[Mux.scala 27:72]
  wire  _T_4908 = btb_rd_addr_p1_f == 8'h55; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5335 = _T_4908 ? _T_985 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5590 = _T_5589 | _T_5335; // @[Mux.scala 27:72]
  wire  _T_4910 = btb_rd_addr_p1_f == 8'h56; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5336 = _T_4910 ? _T_989 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5591 = _T_5590 | _T_5336; // @[Mux.scala 27:72]
  wire  _T_4912 = btb_rd_addr_p1_f == 8'h57; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5337 = _T_4912 ? _T_993 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5592 = _T_5591 | _T_5337; // @[Mux.scala 27:72]
  wire  _T_4914 = btb_rd_addr_p1_f == 8'h58; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5338 = _T_4914 ? _T_997 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5593 = _T_5592 | _T_5338; // @[Mux.scala 27:72]
  wire  _T_4916 = btb_rd_addr_p1_f == 8'h59; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5339 = _T_4916 ? _T_1001 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5594 = _T_5593 | _T_5339; // @[Mux.scala 27:72]
  wire  _T_4918 = btb_rd_addr_p1_f == 8'h5a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5340 = _T_4918 ? _T_1005 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5595 = _T_5594 | _T_5340; // @[Mux.scala 27:72]
  wire  _T_4920 = btb_rd_addr_p1_f == 8'h5b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5341 = _T_4920 ? _T_1009 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5596 = _T_5595 | _T_5341; // @[Mux.scala 27:72]
  wire  _T_4922 = btb_rd_addr_p1_f == 8'h5c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5342 = _T_4922 ? _T_1013 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5597 = _T_5596 | _T_5342; // @[Mux.scala 27:72]
  wire  _T_4924 = btb_rd_addr_p1_f == 8'h5d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5343 = _T_4924 ? _T_1017 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5598 = _T_5597 | _T_5343; // @[Mux.scala 27:72]
  wire  _T_4926 = btb_rd_addr_p1_f == 8'h5e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5344 = _T_4926 ? _T_1021 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5599 = _T_5598 | _T_5344; // @[Mux.scala 27:72]
  wire  _T_4928 = btb_rd_addr_p1_f == 8'h5f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5345 = _T_4928 ? _T_1025 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5600 = _T_5599 | _T_5345; // @[Mux.scala 27:72]
  wire  _T_4930 = btb_rd_addr_p1_f == 8'h60; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5346 = _T_4930 ? _T_1029 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5601 = _T_5600 | _T_5346; // @[Mux.scala 27:72]
  wire  _T_4932 = btb_rd_addr_p1_f == 8'h61; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5347 = _T_4932 ? _T_1033 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5602 = _T_5601 | _T_5347; // @[Mux.scala 27:72]
  wire  _T_4934 = btb_rd_addr_p1_f == 8'h62; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5348 = _T_4934 ? _T_1037 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5603 = _T_5602 | _T_5348; // @[Mux.scala 27:72]
  wire  _T_4936 = btb_rd_addr_p1_f == 8'h63; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5349 = _T_4936 ? _T_1041 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5604 = _T_5603 | _T_5349; // @[Mux.scala 27:72]
  wire  _T_4938 = btb_rd_addr_p1_f == 8'h64; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5350 = _T_4938 ? _T_1045 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5605 = _T_5604 | _T_5350; // @[Mux.scala 27:72]
  wire  _T_4940 = btb_rd_addr_p1_f == 8'h65; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5351 = _T_4940 ? _T_1049 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5606 = _T_5605 | _T_5351; // @[Mux.scala 27:72]
  wire  _T_4942 = btb_rd_addr_p1_f == 8'h66; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5352 = _T_4942 ? _T_1053 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5607 = _T_5606 | _T_5352; // @[Mux.scala 27:72]
  wire  _T_4944 = btb_rd_addr_p1_f == 8'h67; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5353 = _T_4944 ? _T_1057 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5608 = _T_5607 | _T_5353; // @[Mux.scala 27:72]
  wire  _T_4946 = btb_rd_addr_p1_f == 8'h68; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5354 = _T_4946 ? _T_1061 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5609 = _T_5608 | _T_5354; // @[Mux.scala 27:72]
  wire  _T_4948 = btb_rd_addr_p1_f == 8'h69; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5355 = _T_4948 ? _T_1065 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5610 = _T_5609 | _T_5355; // @[Mux.scala 27:72]
  wire  _T_4950 = btb_rd_addr_p1_f == 8'h6a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5356 = _T_4950 ? _T_1069 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5611 = _T_5610 | _T_5356; // @[Mux.scala 27:72]
  wire  _T_4952 = btb_rd_addr_p1_f == 8'h6b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5357 = _T_4952 ? _T_1073 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5612 = _T_5611 | _T_5357; // @[Mux.scala 27:72]
  wire  _T_4954 = btb_rd_addr_p1_f == 8'h6c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5358 = _T_4954 ? _T_1077 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5613 = _T_5612 | _T_5358; // @[Mux.scala 27:72]
  wire  _T_4956 = btb_rd_addr_p1_f == 8'h6d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5359 = _T_4956 ? _T_1081 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5614 = _T_5613 | _T_5359; // @[Mux.scala 27:72]
  wire  _T_4958 = btb_rd_addr_p1_f == 8'h6e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5360 = _T_4958 ? _T_1085 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5615 = _T_5614 | _T_5360; // @[Mux.scala 27:72]
  wire  _T_4960 = btb_rd_addr_p1_f == 8'h6f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5361 = _T_4960 ? _T_1089 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5616 = _T_5615 | _T_5361; // @[Mux.scala 27:72]
  wire  _T_4962 = btb_rd_addr_p1_f == 8'h70; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5362 = _T_4962 ? _T_1093 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5617 = _T_5616 | _T_5362; // @[Mux.scala 27:72]
  wire  _T_4964 = btb_rd_addr_p1_f == 8'h71; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5363 = _T_4964 ? _T_1097 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5618 = _T_5617 | _T_5363; // @[Mux.scala 27:72]
  wire  _T_4966 = btb_rd_addr_p1_f == 8'h72; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5364 = _T_4966 ? _T_1101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5619 = _T_5618 | _T_5364; // @[Mux.scala 27:72]
  wire  _T_4968 = btb_rd_addr_p1_f == 8'h73; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5365 = _T_4968 ? _T_1105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5620 = _T_5619 | _T_5365; // @[Mux.scala 27:72]
  wire  _T_4970 = btb_rd_addr_p1_f == 8'h74; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5366 = _T_4970 ? _T_1109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5621 = _T_5620 | _T_5366; // @[Mux.scala 27:72]
  wire  _T_4972 = btb_rd_addr_p1_f == 8'h75; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5367 = _T_4972 ? _T_1113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5622 = _T_5621 | _T_5367; // @[Mux.scala 27:72]
  wire  _T_4974 = btb_rd_addr_p1_f == 8'h76; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5368 = _T_4974 ? _T_1117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5623 = _T_5622 | _T_5368; // @[Mux.scala 27:72]
  wire  _T_4976 = btb_rd_addr_p1_f == 8'h77; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5369 = _T_4976 ? _T_1121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5624 = _T_5623 | _T_5369; // @[Mux.scala 27:72]
  wire  _T_4978 = btb_rd_addr_p1_f == 8'h78; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5370 = _T_4978 ? _T_1125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5625 = _T_5624 | _T_5370; // @[Mux.scala 27:72]
  wire  _T_4980 = btb_rd_addr_p1_f == 8'h79; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5371 = _T_4980 ? _T_1129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5626 = _T_5625 | _T_5371; // @[Mux.scala 27:72]
  wire  _T_4982 = btb_rd_addr_p1_f == 8'h7a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5372 = _T_4982 ? _T_1133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5627 = _T_5626 | _T_5372; // @[Mux.scala 27:72]
  wire  _T_4984 = btb_rd_addr_p1_f == 8'h7b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5373 = _T_4984 ? _T_1137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5628 = _T_5627 | _T_5373; // @[Mux.scala 27:72]
  wire  _T_4986 = btb_rd_addr_p1_f == 8'h7c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5374 = _T_4986 ? _T_1141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5629 = _T_5628 | _T_5374; // @[Mux.scala 27:72]
  wire  _T_4988 = btb_rd_addr_p1_f == 8'h7d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5375 = _T_4988 ? _T_1145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5630 = _T_5629 | _T_5375; // @[Mux.scala 27:72]
  wire  _T_4990 = btb_rd_addr_p1_f == 8'h7e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5376 = _T_4990 ? _T_1149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5631 = _T_5630 | _T_5376; // @[Mux.scala 27:72]
  wire  _T_4992 = btb_rd_addr_p1_f == 8'h7f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5377 = _T_4992 ? _T_1153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5632 = _T_5631 | _T_5377; // @[Mux.scala 27:72]
  wire  _T_4994 = btb_rd_addr_p1_f == 8'h80; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5378 = _T_4994 ? _T_1157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5633 = _T_5632 | _T_5378; // @[Mux.scala 27:72]
  wire  _T_4996 = btb_rd_addr_p1_f == 8'h81; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5379 = _T_4996 ? _T_1161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5634 = _T_5633 | _T_5379; // @[Mux.scala 27:72]
  wire  _T_4998 = btb_rd_addr_p1_f == 8'h82; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5380 = _T_4998 ? _T_1165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5635 = _T_5634 | _T_5380; // @[Mux.scala 27:72]
  wire  _T_5000 = btb_rd_addr_p1_f == 8'h83; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5381 = _T_5000 ? _T_1169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5636 = _T_5635 | _T_5381; // @[Mux.scala 27:72]
  wire  _T_5002 = btb_rd_addr_p1_f == 8'h84; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5382 = _T_5002 ? _T_1173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5637 = _T_5636 | _T_5382; // @[Mux.scala 27:72]
  wire  _T_5004 = btb_rd_addr_p1_f == 8'h85; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5383 = _T_5004 ? _T_1177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5638 = _T_5637 | _T_5383; // @[Mux.scala 27:72]
  wire  _T_5006 = btb_rd_addr_p1_f == 8'h86; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5384 = _T_5006 ? _T_1181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5639 = _T_5638 | _T_5384; // @[Mux.scala 27:72]
  wire  _T_5008 = btb_rd_addr_p1_f == 8'h87; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5385 = _T_5008 ? _T_1185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5640 = _T_5639 | _T_5385; // @[Mux.scala 27:72]
  wire  _T_5010 = btb_rd_addr_p1_f == 8'h88; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5386 = _T_5010 ? _T_1189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5641 = _T_5640 | _T_5386; // @[Mux.scala 27:72]
  wire  _T_5012 = btb_rd_addr_p1_f == 8'h89; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5387 = _T_5012 ? _T_1193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5642 = _T_5641 | _T_5387; // @[Mux.scala 27:72]
  wire  _T_5014 = btb_rd_addr_p1_f == 8'h8a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5388 = _T_5014 ? _T_1197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5643 = _T_5642 | _T_5388; // @[Mux.scala 27:72]
  wire  _T_5016 = btb_rd_addr_p1_f == 8'h8b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5389 = _T_5016 ? _T_1201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5644 = _T_5643 | _T_5389; // @[Mux.scala 27:72]
  wire  _T_5018 = btb_rd_addr_p1_f == 8'h8c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5390 = _T_5018 ? _T_1205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5645 = _T_5644 | _T_5390; // @[Mux.scala 27:72]
  wire  _T_5020 = btb_rd_addr_p1_f == 8'h8d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5391 = _T_5020 ? _T_1209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5646 = _T_5645 | _T_5391; // @[Mux.scala 27:72]
  wire  _T_5022 = btb_rd_addr_p1_f == 8'h8e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5392 = _T_5022 ? _T_1213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5647 = _T_5646 | _T_5392; // @[Mux.scala 27:72]
  wire  _T_5024 = btb_rd_addr_p1_f == 8'h8f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5393 = _T_5024 ? _T_1217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5648 = _T_5647 | _T_5393; // @[Mux.scala 27:72]
  wire  _T_5026 = btb_rd_addr_p1_f == 8'h90; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5394 = _T_5026 ? _T_1221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5649 = _T_5648 | _T_5394; // @[Mux.scala 27:72]
  wire  _T_5028 = btb_rd_addr_p1_f == 8'h91; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5395 = _T_5028 ? _T_1225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5650 = _T_5649 | _T_5395; // @[Mux.scala 27:72]
  wire  _T_5030 = btb_rd_addr_p1_f == 8'h92; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5396 = _T_5030 ? _T_1229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5651 = _T_5650 | _T_5396; // @[Mux.scala 27:72]
  wire  _T_5032 = btb_rd_addr_p1_f == 8'h93; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5397 = _T_5032 ? _T_1233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5652 = _T_5651 | _T_5397; // @[Mux.scala 27:72]
  wire  _T_5034 = btb_rd_addr_p1_f == 8'h94; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5398 = _T_5034 ? _T_1237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5653 = _T_5652 | _T_5398; // @[Mux.scala 27:72]
  wire  _T_5036 = btb_rd_addr_p1_f == 8'h95; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5399 = _T_5036 ? _T_1241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5654 = _T_5653 | _T_5399; // @[Mux.scala 27:72]
  wire  _T_5038 = btb_rd_addr_p1_f == 8'h96; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5400 = _T_5038 ? _T_1245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5655 = _T_5654 | _T_5400; // @[Mux.scala 27:72]
  wire  _T_5040 = btb_rd_addr_p1_f == 8'h97; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5401 = _T_5040 ? _T_1249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5656 = _T_5655 | _T_5401; // @[Mux.scala 27:72]
  wire  _T_5042 = btb_rd_addr_p1_f == 8'h98; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5402 = _T_5042 ? _T_1253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5657 = _T_5656 | _T_5402; // @[Mux.scala 27:72]
  wire  _T_5044 = btb_rd_addr_p1_f == 8'h99; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5403 = _T_5044 ? _T_1257 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5658 = _T_5657 | _T_5403; // @[Mux.scala 27:72]
  wire  _T_5046 = btb_rd_addr_p1_f == 8'h9a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5404 = _T_5046 ? _T_1261 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5659 = _T_5658 | _T_5404; // @[Mux.scala 27:72]
  wire  _T_5048 = btb_rd_addr_p1_f == 8'h9b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5405 = _T_5048 ? _T_1265 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5660 = _T_5659 | _T_5405; // @[Mux.scala 27:72]
  wire  _T_5050 = btb_rd_addr_p1_f == 8'h9c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5406 = _T_5050 ? _T_1269 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5661 = _T_5660 | _T_5406; // @[Mux.scala 27:72]
  wire  _T_5052 = btb_rd_addr_p1_f == 8'h9d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5407 = _T_5052 ? _T_1273 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5662 = _T_5661 | _T_5407; // @[Mux.scala 27:72]
  wire  _T_5054 = btb_rd_addr_p1_f == 8'h9e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5408 = _T_5054 ? _T_1277 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5663 = _T_5662 | _T_5408; // @[Mux.scala 27:72]
  wire  _T_5056 = btb_rd_addr_p1_f == 8'h9f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5409 = _T_5056 ? _T_1281 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5664 = _T_5663 | _T_5409; // @[Mux.scala 27:72]
  wire  _T_5058 = btb_rd_addr_p1_f == 8'ha0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5410 = _T_5058 ? _T_1285 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5665 = _T_5664 | _T_5410; // @[Mux.scala 27:72]
  wire  _T_5060 = btb_rd_addr_p1_f == 8'ha1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5411 = _T_5060 ? _T_1289 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5666 = _T_5665 | _T_5411; // @[Mux.scala 27:72]
  wire  _T_5062 = btb_rd_addr_p1_f == 8'ha2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5412 = _T_5062 ? _T_1293 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5667 = _T_5666 | _T_5412; // @[Mux.scala 27:72]
  wire  _T_5064 = btb_rd_addr_p1_f == 8'ha3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5413 = _T_5064 ? _T_1297 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5668 = _T_5667 | _T_5413; // @[Mux.scala 27:72]
  wire  _T_5066 = btb_rd_addr_p1_f == 8'ha4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5414 = _T_5066 ? _T_1301 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5669 = _T_5668 | _T_5414; // @[Mux.scala 27:72]
  wire  _T_5068 = btb_rd_addr_p1_f == 8'ha5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5415 = _T_5068 ? _T_1305 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5670 = _T_5669 | _T_5415; // @[Mux.scala 27:72]
  wire  _T_5070 = btb_rd_addr_p1_f == 8'ha6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5416 = _T_5070 ? _T_1309 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5671 = _T_5670 | _T_5416; // @[Mux.scala 27:72]
  wire  _T_5072 = btb_rd_addr_p1_f == 8'ha7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5417 = _T_5072 ? _T_1313 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5672 = _T_5671 | _T_5417; // @[Mux.scala 27:72]
  wire  _T_5074 = btb_rd_addr_p1_f == 8'ha8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5418 = _T_5074 ? _T_1317 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5673 = _T_5672 | _T_5418; // @[Mux.scala 27:72]
  wire  _T_5076 = btb_rd_addr_p1_f == 8'ha9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5419 = _T_5076 ? _T_1321 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5674 = _T_5673 | _T_5419; // @[Mux.scala 27:72]
  wire  _T_5078 = btb_rd_addr_p1_f == 8'haa; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5420 = _T_5078 ? _T_1325 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5675 = _T_5674 | _T_5420; // @[Mux.scala 27:72]
  wire  _T_5080 = btb_rd_addr_p1_f == 8'hab; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5421 = _T_5080 ? _T_1329 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5676 = _T_5675 | _T_5421; // @[Mux.scala 27:72]
  wire  _T_5082 = btb_rd_addr_p1_f == 8'hac; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5422 = _T_5082 ? _T_1333 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5677 = _T_5676 | _T_5422; // @[Mux.scala 27:72]
  wire  _T_5084 = btb_rd_addr_p1_f == 8'had; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5423 = _T_5084 ? _T_1337 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5678 = _T_5677 | _T_5423; // @[Mux.scala 27:72]
  wire  _T_5086 = btb_rd_addr_p1_f == 8'hae; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5424 = _T_5086 ? _T_1341 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5679 = _T_5678 | _T_5424; // @[Mux.scala 27:72]
  wire  _T_5088 = btb_rd_addr_p1_f == 8'haf; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5425 = _T_5088 ? _T_1345 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5680 = _T_5679 | _T_5425; // @[Mux.scala 27:72]
  wire  _T_5090 = btb_rd_addr_p1_f == 8'hb0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5426 = _T_5090 ? _T_1349 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5681 = _T_5680 | _T_5426; // @[Mux.scala 27:72]
  wire  _T_5092 = btb_rd_addr_p1_f == 8'hb1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5427 = _T_5092 ? _T_1353 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5682 = _T_5681 | _T_5427; // @[Mux.scala 27:72]
  wire  _T_5094 = btb_rd_addr_p1_f == 8'hb2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5428 = _T_5094 ? _T_1357 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5683 = _T_5682 | _T_5428; // @[Mux.scala 27:72]
  wire  _T_5096 = btb_rd_addr_p1_f == 8'hb3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5429 = _T_5096 ? _T_1361 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5684 = _T_5683 | _T_5429; // @[Mux.scala 27:72]
  wire  _T_5098 = btb_rd_addr_p1_f == 8'hb4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5430 = _T_5098 ? _T_1365 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5685 = _T_5684 | _T_5430; // @[Mux.scala 27:72]
  wire  _T_5100 = btb_rd_addr_p1_f == 8'hb5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5431 = _T_5100 ? _T_1369 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5686 = _T_5685 | _T_5431; // @[Mux.scala 27:72]
  wire  _T_5102 = btb_rd_addr_p1_f == 8'hb6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5432 = _T_5102 ? _T_1373 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5687 = _T_5686 | _T_5432; // @[Mux.scala 27:72]
  wire  _T_5104 = btb_rd_addr_p1_f == 8'hb7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5433 = _T_5104 ? _T_1377 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5688 = _T_5687 | _T_5433; // @[Mux.scala 27:72]
  wire  _T_5106 = btb_rd_addr_p1_f == 8'hb8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5434 = _T_5106 ? _T_1381 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5689 = _T_5688 | _T_5434; // @[Mux.scala 27:72]
  wire  _T_5108 = btb_rd_addr_p1_f == 8'hb9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5435 = _T_5108 ? _T_1385 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5690 = _T_5689 | _T_5435; // @[Mux.scala 27:72]
  wire  _T_5110 = btb_rd_addr_p1_f == 8'hba; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5436 = _T_5110 ? _T_1389 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5691 = _T_5690 | _T_5436; // @[Mux.scala 27:72]
  wire  _T_5112 = btb_rd_addr_p1_f == 8'hbb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5437 = _T_5112 ? _T_1393 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5692 = _T_5691 | _T_5437; // @[Mux.scala 27:72]
  wire  _T_5114 = btb_rd_addr_p1_f == 8'hbc; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5438 = _T_5114 ? _T_1397 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5693 = _T_5692 | _T_5438; // @[Mux.scala 27:72]
  wire  _T_5116 = btb_rd_addr_p1_f == 8'hbd; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5439 = _T_5116 ? _T_1401 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5694 = _T_5693 | _T_5439; // @[Mux.scala 27:72]
  wire  _T_5118 = btb_rd_addr_p1_f == 8'hbe; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5440 = _T_5118 ? _T_1405 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5695 = _T_5694 | _T_5440; // @[Mux.scala 27:72]
  wire  _T_5120 = btb_rd_addr_p1_f == 8'hbf; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5441 = _T_5120 ? _T_1409 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5696 = _T_5695 | _T_5441; // @[Mux.scala 27:72]
  wire  _T_5122 = btb_rd_addr_p1_f == 8'hc0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5442 = _T_5122 ? _T_1413 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5697 = _T_5696 | _T_5442; // @[Mux.scala 27:72]
  wire  _T_5124 = btb_rd_addr_p1_f == 8'hc1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5443 = _T_5124 ? _T_1417 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5698 = _T_5697 | _T_5443; // @[Mux.scala 27:72]
  wire  _T_5126 = btb_rd_addr_p1_f == 8'hc2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5444 = _T_5126 ? _T_1421 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5699 = _T_5698 | _T_5444; // @[Mux.scala 27:72]
  wire  _T_5128 = btb_rd_addr_p1_f == 8'hc3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5445 = _T_5128 ? _T_1425 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5700 = _T_5699 | _T_5445; // @[Mux.scala 27:72]
  wire  _T_5130 = btb_rd_addr_p1_f == 8'hc4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5446 = _T_5130 ? _T_1429 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5701 = _T_5700 | _T_5446; // @[Mux.scala 27:72]
  wire  _T_5132 = btb_rd_addr_p1_f == 8'hc5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5447 = _T_5132 ? _T_1433 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5702 = _T_5701 | _T_5447; // @[Mux.scala 27:72]
  wire  _T_5134 = btb_rd_addr_p1_f == 8'hc6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5448 = _T_5134 ? _T_1437 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5703 = _T_5702 | _T_5448; // @[Mux.scala 27:72]
  wire  _T_5136 = btb_rd_addr_p1_f == 8'hc7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5449 = _T_5136 ? _T_1441 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5704 = _T_5703 | _T_5449; // @[Mux.scala 27:72]
  wire  _T_5138 = btb_rd_addr_p1_f == 8'hc8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5450 = _T_5138 ? _T_1445 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5705 = _T_5704 | _T_5450; // @[Mux.scala 27:72]
  wire  _T_5140 = btb_rd_addr_p1_f == 8'hc9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5451 = _T_5140 ? _T_1449 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5706 = _T_5705 | _T_5451; // @[Mux.scala 27:72]
  wire  _T_5142 = btb_rd_addr_p1_f == 8'hca; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5452 = _T_5142 ? _T_1453 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5707 = _T_5706 | _T_5452; // @[Mux.scala 27:72]
  wire  _T_5144 = btb_rd_addr_p1_f == 8'hcb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5453 = _T_5144 ? _T_1457 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5708 = _T_5707 | _T_5453; // @[Mux.scala 27:72]
  wire  _T_5146 = btb_rd_addr_p1_f == 8'hcc; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5454 = _T_5146 ? _T_1461 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5709 = _T_5708 | _T_5454; // @[Mux.scala 27:72]
  wire  _T_5148 = btb_rd_addr_p1_f == 8'hcd; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5455 = _T_5148 ? _T_1465 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5710 = _T_5709 | _T_5455; // @[Mux.scala 27:72]
  wire  _T_5150 = btb_rd_addr_p1_f == 8'hce; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5456 = _T_5150 ? _T_1469 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5711 = _T_5710 | _T_5456; // @[Mux.scala 27:72]
  wire  _T_5152 = btb_rd_addr_p1_f == 8'hcf; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5457 = _T_5152 ? _T_1473 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5712 = _T_5711 | _T_5457; // @[Mux.scala 27:72]
  wire  _T_5154 = btb_rd_addr_p1_f == 8'hd0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5458 = _T_5154 ? _T_1477 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5713 = _T_5712 | _T_5458; // @[Mux.scala 27:72]
  wire  _T_5156 = btb_rd_addr_p1_f == 8'hd1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5459 = _T_5156 ? _T_1481 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5714 = _T_5713 | _T_5459; // @[Mux.scala 27:72]
  wire  _T_5158 = btb_rd_addr_p1_f == 8'hd2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5460 = _T_5158 ? _T_1485 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5715 = _T_5714 | _T_5460; // @[Mux.scala 27:72]
  wire  _T_5160 = btb_rd_addr_p1_f == 8'hd3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5461 = _T_5160 ? _T_1489 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5716 = _T_5715 | _T_5461; // @[Mux.scala 27:72]
  wire  _T_5162 = btb_rd_addr_p1_f == 8'hd4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5462 = _T_5162 ? _T_1493 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5717 = _T_5716 | _T_5462; // @[Mux.scala 27:72]
  wire  _T_5164 = btb_rd_addr_p1_f == 8'hd5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5463 = _T_5164 ? _T_1497 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5718 = _T_5717 | _T_5463; // @[Mux.scala 27:72]
  wire  _T_5166 = btb_rd_addr_p1_f == 8'hd6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5464 = _T_5166 ? _T_1501 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5719 = _T_5718 | _T_5464; // @[Mux.scala 27:72]
  wire  _T_5168 = btb_rd_addr_p1_f == 8'hd7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5465 = _T_5168 ? _T_1505 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5720 = _T_5719 | _T_5465; // @[Mux.scala 27:72]
  wire  _T_5170 = btb_rd_addr_p1_f == 8'hd8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5466 = _T_5170 ? _T_1509 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5721 = _T_5720 | _T_5466; // @[Mux.scala 27:72]
  wire  _T_5172 = btb_rd_addr_p1_f == 8'hd9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5467 = _T_5172 ? _T_1513 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5722 = _T_5721 | _T_5467; // @[Mux.scala 27:72]
  wire  _T_5174 = btb_rd_addr_p1_f == 8'hda; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5468 = _T_5174 ? _T_1517 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5723 = _T_5722 | _T_5468; // @[Mux.scala 27:72]
  wire  _T_5176 = btb_rd_addr_p1_f == 8'hdb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5469 = _T_5176 ? _T_1521 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5724 = _T_5723 | _T_5469; // @[Mux.scala 27:72]
  wire  _T_5178 = btb_rd_addr_p1_f == 8'hdc; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5470 = _T_5178 ? _T_1525 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5725 = _T_5724 | _T_5470; // @[Mux.scala 27:72]
  wire  _T_5180 = btb_rd_addr_p1_f == 8'hdd; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5471 = _T_5180 ? _T_1529 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5726 = _T_5725 | _T_5471; // @[Mux.scala 27:72]
  wire  _T_5182 = btb_rd_addr_p1_f == 8'hde; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5472 = _T_5182 ? _T_1533 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5727 = _T_5726 | _T_5472; // @[Mux.scala 27:72]
  wire  _T_5184 = btb_rd_addr_p1_f == 8'hdf; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5473 = _T_5184 ? _T_1537 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5728 = _T_5727 | _T_5473; // @[Mux.scala 27:72]
  wire  _T_5186 = btb_rd_addr_p1_f == 8'he0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5474 = _T_5186 ? _T_1541 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5729 = _T_5728 | _T_5474; // @[Mux.scala 27:72]
  wire  _T_5188 = btb_rd_addr_p1_f == 8'he1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5475 = _T_5188 ? _T_1545 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5730 = _T_5729 | _T_5475; // @[Mux.scala 27:72]
  wire  _T_5190 = btb_rd_addr_p1_f == 8'he2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5476 = _T_5190 ? _T_1549 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5731 = _T_5730 | _T_5476; // @[Mux.scala 27:72]
  wire  _T_5192 = btb_rd_addr_p1_f == 8'he3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5477 = _T_5192 ? _T_1553 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5732 = _T_5731 | _T_5477; // @[Mux.scala 27:72]
  wire  _T_5194 = btb_rd_addr_p1_f == 8'he4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5478 = _T_5194 ? _T_1557 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5733 = _T_5732 | _T_5478; // @[Mux.scala 27:72]
  wire  _T_5196 = btb_rd_addr_p1_f == 8'he5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5479 = _T_5196 ? _T_1561 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5734 = _T_5733 | _T_5479; // @[Mux.scala 27:72]
  wire  _T_5198 = btb_rd_addr_p1_f == 8'he6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5480 = _T_5198 ? _T_1565 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5735 = _T_5734 | _T_5480; // @[Mux.scala 27:72]
  wire  _T_5200 = btb_rd_addr_p1_f == 8'he7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5481 = _T_5200 ? _T_1569 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5736 = _T_5735 | _T_5481; // @[Mux.scala 27:72]
  wire  _T_5202 = btb_rd_addr_p1_f == 8'he8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5482 = _T_5202 ? _T_1573 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5737 = _T_5736 | _T_5482; // @[Mux.scala 27:72]
  wire  _T_5204 = btb_rd_addr_p1_f == 8'he9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5483 = _T_5204 ? _T_1577 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5738 = _T_5737 | _T_5483; // @[Mux.scala 27:72]
  wire  _T_5206 = btb_rd_addr_p1_f == 8'hea; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5484 = _T_5206 ? _T_1581 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5739 = _T_5738 | _T_5484; // @[Mux.scala 27:72]
  wire  _T_5208 = btb_rd_addr_p1_f == 8'heb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5485 = _T_5208 ? _T_1585 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5740 = _T_5739 | _T_5485; // @[Mux.scala 27:72]
  wire  _T_5210 = btb_rd_addr_p1_f == 8'hec; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5486 = _T_5210 ? _T_1589 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5741 = _T_5740 | _T_5486; // @[Mux.scala 27:72]
  wire  _T_5212 = btb_rd_addr_p1_f == 8'hed; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5487 = _T_5212 ? _T_1593 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5742 = _T_5741 | _T_5487; // @[Mux.scala 27:72]
  wire  _T_5214 = btb_rd_addr_p1_f == 8'hee; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5488 = _T_5214 ? _T_1597 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5743 = _T_5742 | _T_5488; // @[Mux.scala 27:72]
  wire  _T_5216 = btb_rd_addr_p1_f == 8'hef; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5489 = _T_5216 ? _T_1601 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5744 = _T_5743 | _T_5489; // @[Mux.scala 27:72]
  wire  _T_5218 = btb_rd_addr_p1_f == 8'hf0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5490 = _T_5218 ? _T_1605 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5745 = _T_5744 | _T_5490; // @[Mux.scala 27:72]
  wire  _T_5220 = btb_rd_addr_p1_f == 8'hf1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5491 = _T_5220 ? _T_1609 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5746 = _T_5745 | _T_5491; // @[Mux.scala 27:72]
  wire  _T_5222 = btb_rd_addr_p1_f == 8'hf2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5492 = _T_5222 ? _T_1613 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5747 = _T_5746 | _T_5492; // @[Mux.scala 27:72]
  wire  _T_5224 = btb_rd_addr_p1_f == 8'hf3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5493 = _T_5224 ? _T_1617 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5748 = _T_5747 | _T_5493; // @[Mux.scala 27:72]
  wire  _T_5226 = btb_rd_addr_p1_f == 8'hf4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5494 = _T_5226 ? _T_1621 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5749 = _T_5748 | _T_5494; // @[Mux.scala 27:72]
  wire  _T_5228 = btb_rd_addr_p1_f == 8'hf5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5495 = _T_5228 ? _T_1625 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5750 = _T_5749 | _T_5495; // @[Mux.scala 27:72]
  wire  _T_5230 = btb_rd_addr_p1_f == 8'hf6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5496 = _T_5230 ? _T_1629 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5751 = _T_5750 | _T_5496; // @[Mux.scala 27:72]
  wire  _T_5232 = btb_rd_addr_p1_f == 8'hf7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5497 = _T_5232 ? _T_1633 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5752 = _T_5751 | _T_5497; // @[Mux.scala 27:72]
  wire  _T_5234 = btb_rd_addr_p1_f == 8'hf8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5498 = _T_5234 ? _T_1637 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5753 = _T_5752 | _T_5498; // @[Mux.scala 27:72]
  wire  _T_5236 = btb_rd_addr_p1_f == 8'hf9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5499 = _T_5236 ? _T_1641 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5754 = _T_5753 | _T_5499; // @[Mux.scala 27:72]
  wire  _T_5238 = btb_rd_addr_p1_f == 8'hfa; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5500 = _T_5238 ? _T_1645 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5755 = _T_5754 | _T_5500; // @[Mux.scala 27:72]
  wire  _T_5240 = btb_rd_addr_p1_f == 8'hfb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5501 = _T_5240 ? _T_1649 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5756 = _T_5755 | _T_5501; // @[Mux.scala 27:72]
  wire  _T_5242 = btb_rd_addr_p1_f == 8'hfc; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5502 = _T_5242 ? _T_1653 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5757 = _T_5756 | _T_5502; // @[Mux.scala 27:72]
  wire  _T_5244 = btb_rd_addr_p1_f == 8'hfd; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5503 = _T_5244 ? _T_1657 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5758 = _T_5757 | _T_5503; // @[Mux.scala 27:72]
  wire  _T_5246 = btb_rd_addr_p1_f == 8'hfe; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5504 = _T_5246 ? _T_1661 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5759 = _T_5758 | _T_5504; // @[Mux.scala 27:72]
  wire  _T_5248 = btb_rd_addr_p1_f == 8'hff; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_5505 = _T_5248 ? _T_1665 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5760 = _T_5759 | _T_5505; // @[Mux.scala 27:72]
  wire [21:0] _T_5761 = _T_5760; // @[Mux.scala 27:72 Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_p1_f = _T_5760; // @[ifu_bp_ctl.scala 441:31]
  wire [4:0] _T_36 = _T_8[13:9] ^ _T_8[18:14]; // @[lib.scala 42:111]
  wire [4:0] _T_37 = _T_36 ^ _T_8[23:19]; // @[lib.scala 42:111]
  wire  _T_70 = _T_5761[21:17] == _T_37; // @[ifu_bp_ctl.scala 152:107]
  wire  _T_71 = _T_5761[0] & _T_70; // @[ifu_bp_ctl.scala 152:61]
  wire  _T_20 = io_exu_bp_exu_i0_br_index_r == btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 126:75]
  wire  branch_error_collision_p1_f = dec_tlu_error_wb & _T_20; // @[ifu_bp_ctl.scala 126:54]
  wire  branch_error_bank_conflict_p1_f = branch_error_collision_p1_f & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 130:69]
  wire  _T_72 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & branch_error_bank_conflict_p1_f; // @[ifu_bp_ctl.scala 153:22]
  wire  _T_73 = ~_T_72; // @[ifu_bp_ctl.scala 153:5]
  wire  _T_74 = _T_71 & _T_73; // @[ifu_bp_ctl.scala 152:130]
  wire  _T_75 = _T_74 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 153:57]
  wire  _T_77 = _T_75 & _T; // @[ifu_bp_ctl.scala 153:78]
  wire  _T_110 = _T_5761[3] ^ _T_5761[4]; // @[ifu_bp_ctl.scala 165:99]
  wire  _T_111 = _T_77 & _T_110; // @[ifu_bp_ctl.scala 165:62]
  wire  _T_115 = ~_T_110; // @[ifu_bp_ctl.scala 166:27]
  wire  _T_116 = _T_77 & _T_115; // @[ifu_bp_ctl.scala 166:25]
  wire [1:0] _T_117 = {_T_111,_T_116}; // @[Cat.scala 29:58]
  wire [21:0] _T_150 = _T_117[0] ? _T_5761 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6274 = _T_4738 ? _T_1669 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6275 = _T_4740 ? _T_1673 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6530 = _T_6274 | _T_6275; // @[Mux.scala 27:72]
  wire [21:0] _T_6276 = _T_4742 ? _T_1677 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6531 = _T_6530 | _T_6276; // @[Mux.scala 27:72]
  wire [21:0] _T_6277 = _T_4744 ? _T_1681 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6532 = _T_6531 | _T_6277; // @[Mux.scala 27:72]
  wire [21:0] _T_6278 = _T_4746 ? _T_1685 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6533 = _T_6532 | _T_6278; // @[Mux.scala 27:72]
  wire [21:0] _T_6279 = _T_4748 ? _T_1689 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6534 = _T_6533 | _T_6279; // @[Mux.scala 27:72]
  wire [21:0] _T_6280 = _T_4750 ? _T_1693 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6535 = _T_6534 | _T_6280; // @[Mux.scala 27:72]
  wire [21:0] _T_6281 = _T_4752 ? _T_1697 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6536 = _T_6535 | _T_6281; // @[Mux.scala 27:72]
  wire [21:0] _T_6282 = _T_4754 ? _T_1701 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6537 = _T_6536 | _T_6282; // @[Mux.scala 27:72]
  wire [21:0] _T_6283 = _T_4756 ? _T_1705 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6538 = _T_6537 | _T_6283; // @[Mux.scala 27:72]
  wire [21:0] _T_6284 = _T_4758 ? _T_1709 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6539 = _T_6538 | _T_6284; // @[Mux.scala 27:72]
  wire [21:0] _T_6285 = _T_4760 ? _T_1713 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6540 = _T_6539 | _T_6285; // @[Mux.scala 27:72]
  wire [21:0] _T_6286 = _T_4762 ? _T_1717 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6541 = _T_6540 | _T_6286; // @[Mux.scala 27:72]
  wire [21:0] _T_6287 = _T_4764 ? _T_1721 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6542 = _T_6541 | _T_6287; // @[Mux.scala 27:72]
  wire [21:0] _T_6288 = _T_4766 ? _T_1725 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6543 = _T_6542 | _T_6288; // @[Mux.scala 27:72]
  wire [21:0] _T_6289 = _T_4768 ? _T_1729 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6544 = _T_6543 | _T_6289; // @[Mux.scala 27:72]
  wire [21:0] _T_6290 = _T_4770 ? _T_1733 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6545 = _T_6544 | _T_6290; // @[Mux.scala 27:72]
  wire [21:0] _T_6291 = _T_4772 ? _T_1737 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6546 = _T_6545 | _T_6291; // @[Mux.scala 27:72]
  wire [21:0] _T_6292 = _T_4774 ? _T_1741 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6547 = _T_6546 | _T_6292; // @[Mux.scala 27:72]
  wire [21:0] _T_6293 = _T_4776 ? _T_1745 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6548 = _T_6547 | _T_6293; // @[Mux.scala 27:72]
  wire [21:0] _T_6294 = _T_4778 ? _T_1749 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6549 = _T_6548 | _T_6294; // @[Mux.scala 27:72]
  wire [21:0] _T_6295 = _T_4780 ? _T_1753 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6550 = _T_6549 | _T_6295; // @[Mux.scala 27:72]
  wire [21:0] _T_6296 = _T_4782 ? _T_1757 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6551 = _T_6550 | _T_6296; // @[Mux.scala 27:72]
  wire [21:0] _T_6297 = _T_4784 ? _T_1761 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6552 = _T_6551 | _T_6297; // @[Mux.scala 27:72]
  wire [21:0] _T_6298 = _T_4786 ? _T_1765 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6553 = _T_6552 | _T_6298; // @[Mux.scala 27:72]
  wire [21:0] _T_6299 = _T_4788 ? _T_1769 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6554 = _T_6553 | _T_6299; // @[Mux.scala 27:72]
  wire [21:0] _T_6300 = _T_4790 ? _T_1773 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6555 = _T_6554 | _T_6300; // @[Mux.scala 27:72]
  wire [21:0] _T_6301 = _T_4792 ? _T_1777 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6556 = _T_6555 | _T_6301; // @[Mux.scala 27:72]
  wire [21:0] _T_6302 = _T_4794 ? _T_1781 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6557 = _T_6556 | _T_6302; // @[Mux.scala 27:72]
  wire [21:0] _T_6303 = _T_4796 ? _T_1785 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6558 = _T_6557 | _T_6303; // @[Mux.scala 27:72]
  wire [21:0] _T_6304 = _T_4798 ? _T_1789 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6559 = _T_6558 | _T_6304; // @[Mux.scala 27:72]
  wire [21:0] _T_6305 = _T_4800 ? _T_1793 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6560 = _T_6559 | _T_6305; // @[Mux.scala 27:72]
  wire [21:0] _T_6306 = _T_4802 ? _T_1797 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6561 = _T_6560 | _T_6306; // @[Mux.scala 27:72]
  wire [21:0] _T_6307 = _T_4804 ? _T_1801 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6562 = _T_6561 | _T_6307; // @[Mux.scala 27:72]
  wire [21:0] _T_6308 = _T_4806 ? _T_1805 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6563 = _T_6562 | _T_6308; // @[Mux.scala 27:72]
  wire [21:0] _T_6309 = _T_4808 ? _T_1809 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6564 = _T_6563 | _T_6309; // @[Mux.scala 27:72]
  wire [21:0] _T_6310 = _T_4810 ? _T_1813 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6565 = _T_6564 | _T_6310; // @[Mux.scala 27:72]
  wire [21:0] _T_6311 = _T_4812 ? _T_1817 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6566 = _T_6565 | _T_6311; // @[Mux.scala 27:72]
  wire [21:0] _T_6312 = _T_4814 ? _T_1821 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6567 = _T_6566 | _T_6312; // @[Mux.scala 27:72]
  wire [21:0] _T_6313 = _T_4816 ? _T_1825 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6568 = _T_6567 | _T_6313; // @[Mux.scala 27:72]
  wire [21:0] _T_6314 = _T_4818 ? _T_1829 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6569 = _T_6568 | _T_6314; // @[Mux.scala 27:72]
  wire [21:0] _T_6315 = _T_4820 ? _T_1833 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6570 = _T_6569 | _T_6315; // @[Mux.scala 27:72]
  wire [21:0] _T_6316 = _T_4822 ? _T_1837 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6571 = _T_6570 | _T_6316; // @[Mux.scala 27:72]
  wire [21:0] _T_6317 = _T_4824 ? _T_1841 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6572 = _T_6571 | _T_6317; // @[Mux.scala 27:72]
  wire [21:0] _T_6318 = _T_4826 ? _T_1845 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6573 = _T_6572 | _T_6318; // @[Mux.scala 27:72]
  wire [21:0] _T_6319 = _T_4828 ? _T_1849 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6574 = _T_6573 | _T_6319; // @[Mux.scala 27:72]
  wire [21:0] _T_6320 = _T_4830 ? _T_1853 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6575 = _T_6574 | _T_6320; // @[Mux.scala 27:72]
  wire [21:0] _T_6321 = _T_4832 ? _T_1857 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6576 = _T_6575 | _T_6321; // @[Mux.scala 27:72]
  wire [21:0] _T_6322 = _T_4834 ? _T_1861 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6577 = _T_6576 | _T_6322; // @[Mux.scala 27:72]
  wire [21:0] _T_6323 = _T_4836 ? _T_1865 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6578 = _T_6577 | _T_6323; // @[Mux.scala 27:72]
  wire [21:0] _T_6324 = _T_4838 ? _T_1869 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6579 = _T_6578 | _T_6324; // @[Mux.scala 27:72]
  wire [21:0] _T_6325 = _T_4840 ? _T_1873 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6580 = _T_6579 | _T_6325; // @[Mux.scala 27:72]
  wire [21:0] _T_6326 = _T_4842 ? _T_1877 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6581 = _T_6580 | _T_6326; // @[Mux.scala 27:72]
  wire [21:0] _T_6327 = _T_4844 ? _T_1881 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6582 = _T_6581 | _T_6327; // @[Mux.scala 27:72]
  wire [21:0] _T_6328 = _T_4846 ? _T_1885 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6583 = _T_6582 | _T_6328; // @[Mux.scala 27:72]
  wire [21:0] _T_6329 = _T_4848 ? _T_1889 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6584 = _T_6583 | _T_6329; // @[Mux.scala 27:72]
  wire [21:0] _T_6330 = _T_4850 ? _T_1893 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6585 = _T_6584 | _T_6330; // @[Mux.scala 27:72]
  wire [21:0] _T_6331 = _T_4852 ? _T_1897 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6586 = _T_6585 | _T_6331; // @[Mux.scala 27:72]
  wire [21:0] _T_6332 = _T_4854 ? _T_1901 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6587 = _T_6586 | _T_6332; // @[Mux.scala 27:72]
  wire [21:0] _T_6333 = _T_4856 ? _T_1905 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6588 = _T_6587 | _T_6333; // @[Mux.scala 27:72]
  wire [21:0] _T_6334 = _T_4858 ? _T_1909 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6589 = _T_6588 | _T_6334; // @[Mux.scala 27:72]
  wire [21:0] _T_6335 = _T_4860 ? _T_1913 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6590 = _T_6589 | _T_6335; // @[Mux.scala 27:72]
  wire [21:0] _T_6336 = _T_4862 ? _T_1917 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6591 = _T_6590 | _T_6336; // @[Mux.scala 27:72]
  wire [21:0] _T_6337 = _T_4864 ? _T_1921 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6592 = _T_6591 | _T_6337; // @[Mux.scala 27:72]
  wire [21:0] _T_6338 = _T_4866 ? _T_1925 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6593 = _T_6592 | _T_6338; // @[Mux.scala 27:72]
  wire [21:0] _T_6339 = _T_4868 ? _T_1929 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6594 = _T_6593 | _T_6339; // @[Mux.scala 27:72]
  wire [21:0] _T_6340 = _T_4870 ? _T_1933 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6595 = _T_6594 | _T_6340; // @[Mux.scala 27:72]
  wire [21:0] _T_6341 = _T_4872 ? _T_1937 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6596 = _T_6595 | _T_6341; // @[Mux.scala 27:72]
  wire [21:0] _T_6342 = _T_4874 ? _T_1941 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6597 = _T_6596 | _T_6342; // @[Mux.scala 27:72]
  wire [21:0] _T_6343 = _T_4876 ? _T_1945 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6598 = _T_6597 | _T_6343; // @[Mux.scala 27:72]
  wire [21:0] _T_6344 = _T_4878 ? _T_1949 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6599 = _T_6598 | _T_6344; // @[Mux.scala 27:72]
  wire [21:0] _T_6345 = _T_4880 ? _T_1953 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6600 = _T_6599 | _T_6345; // @[Mux.scala 27:72]
  wire [21:0] _T_6346 = _T_4882 ? _T_1957 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6601 = _T_6600 | _T_6346; // @[Mux.scala 27:72]
  wire [21:0] _T_6347 = _T_4884 ? _T_1961 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6602 = _T_6601 | _T_6347; // @[Mux.scala 27:72]
  wire [21:0] _T_6348 = _T_4886 ? _T_1965 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6603 = _T_6602 | _T_6348; // @[Mux.scala 27:72]
  wire [21:0] _T_6349 = _T_4888 ? _T_1969 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6604 = _T_6603 | _T_6349; // @[Mux.scala 27:72]
  wire [21:0] _T_6350 = _T_4890 ? _T_1973 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6605 = _T_6604 | _T_6350; // @[Mux.scala 27:72]
  wire [21:0] _T_6351 = _T_4892 ? _T_1977 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6606 = _T_6605 | _T_6351; // @[Mux.scala 27:72]
  wire [21:0] _T_6352 = _T_4894 ? _T_1981 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6607 = _T_6606 | _T_6352; // @[Mux.scala 27:72]
  wire [21:0] _T_6353 = _T_4896 ? _T_1985 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6608 = _T_6607 | _T_6353; // @[Mux.scala 27:72]
  wire [21:0] _T_6354 = _T_4898 ? _T_1989 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6609 = _T_6608 | _T_6354; // @[Mux.scala 27:72]
  wire [21:0] _T_6355 = _T_4900 ? _T_1993 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6610 = _T_6609 | _T_6355; // @[Mux.scala 27:72]
  wire [21:0] _T_6356 = _T_4902 ? _T_1997 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6611 = _T_6610 | _T_6356; // @[Mux.scala 27:72]
  wire [21:0] _T_6357 = _T_4904 ? _T_2001 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6612 = _T_6611 | _T_6357; // @[Mux.scala 27:72]
  wire [21:0] _T_6358 = _T_4906 ? _T_2005 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6613 = _T_6612 | _T_6358; // @[Mux.scala 27:72]
  wire [21:0] _T_6359 = _T_4908 ? _T_2009 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6614 = _T_6613 | _T_6359; // @[Mux.scala 27:72]
  wire [21:0] _T_6360 = _T_4910 ? _T_2013 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6615 = _T_6614 | _T_6360; // @[Mux.scala 27:72]
  wire [21:0] _T_6361 = _T_4912 ? _T_2017 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6616 = _T_6615 | _T_6361; // @[Mux.scala 27:72]
  wire [21:0] _T_6362 = _T_4914 ? _T_2021 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6617 = _T_6616 | _T_6362; // @[Mux.scala 27:72]
  wire [21:0] _T_6363 = _T_4916 ? _T_2025 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6618 = _T_6617 | _T_6363; // @[Mux.scala 27:72]
  wire [21:0] _T_6364 = _T_4918 ? _T_2029 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6619 = _T_6618 | _T_6364; // @[Mux.scala 27:72]
  wire [21:0] _T_6365 = _T_4920 ? _T_2033 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6620 = _T_6619 | _T_6365; // @[Mux.scala 27:72]
  wire [21:0] _T_6366 = _T_4922 ? _T_2037 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6621 = _T_6620 | _T_6366; // @[Mux.scala 27:72]
  wire [21:0] _T_6367 = _T_4924 ? _T_2041 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6622 = _T_6621 | _T_6367; // @[Mux.scala 27:72]
  wire [21:0] _T_6368 = _T_4926 ? _T_2045 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6623 = _T_6622 | _T_6368; // @[Mux.scala 27:72]
  wire [21:0] _T_6369 = _T_4928 ? _T_2049 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6624 = _T_6623 | _T_6369; // @[Mux.scala 27:72]
  wire [21:0] _T_6370 = _T_4930 ? _T_2053 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6625 = _T_6624 | _T_6370; // @[Mux.scala 27:72]
  wire [21:0] _T_6371 = _T_4932 ? _T_2057 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6626 = _T_6625 | _T_6371; // @[Mux.scala 27:72]
  wire [21:0] _T_6372 = _T_4934 ? _T_2061 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6627 = _T_6626 | _T_6372; // @[Mux.scala 27:72]
  wire [21:0] _T_6373 = _T_4936 ? _T_2065 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6628 = _T_6627 | _T_6373; // @[Mux.scala 27:72]
  wire [21:0] _T_6374 = _T_4938 ? _T_2069 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6629 = _T_6628 | _T_6374; // @[Mux.scala 27:72]
  wire [21:0] _T_6375 = _T_4940 ? _T_2073 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6630 = _T_6629 | _T_6375; // @[Mux.scala 27:72]
  wire [21:0] _T_6376 = _T_4942 ? _T_2077 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6631 = _T_6630 | _T_6376; // @[Mux.scala 27:72]
  wire [21:0] _T_6377 = _T_4944 ? _T_2081 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6632 = _T_6631 | _T_6377; // @[Mux.scala 27:72]
  wire [21:0] _T_6378 = _T_4946 ? _T_2085 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6633 = _T_6632 | _T_6378; // @[Mux.scala 27:72]
  wire [21:0] _T_6379 = _T_4948 ? _T_2089 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6634 = _T_6633 | _T_6379; // @[Mux.scala 27:72]
  wire [21:0] _T_6380 = _T_4950 ? _T_2093 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6635 = _T_6634 | _T_6380; // @[Mux.scala 27:72]
  wire [21:0] _T_6381 = _T_4952 ? _T_2097 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6636 = _T_6635 | _T_6381; // @[Mux.scala 27:72]
  wire [21:0] _T_6382 = _T_4954 ? _T_2101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6637 = _T_6636 | _T_6382; // @[Mux.scala 27:72]
  wire [21:0] _T_6383 = _T_4956 ? _T_2105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6638 = _T_6637 | _T_6383; // @[Mux.scala 27:72]
  wire [21:0] _T_6384 = _T_4958 ? _T_2109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6639 = _T_6638 | _T_6384; // @[Mux.scala 27:72]
  wire [21:0] _T_6385 = _T_4960 ? _T_2113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6640 = _T_6639 | _T_6385; // @[Mux.scala 27:72]
  wire [21:0] _T_6386 = _T_4962 ? _T_2117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6641 = _T_6640 | _T_6386; // @[Mux.scala 27:72]
  wire [21:0] _T_6387 = _T_4964 ? _T_2121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6642 = _T_6641 | _T_6387; // @[Mux.scala 27:72]
  wire [21:0] _T_6388 = _T_4966 ? _T_2125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6643 = _T_6642 | _T_6388; // @[Mux.scala 27:72]
  wire [21:0] _T_6389 = _T_4968 ? _T_2129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6644 = _T_6643 | _T_6389; // @[Mux.scala 27:72]
  wire [21:0] _T_6390 = _T_4970 ? _T_2133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6645 = _T_6644 | _T_6390; // @[Mux.scala 27:72]
  wire [21:0] _T_6391 = _T_4972 ? _T_2137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6646 = _T_6645 | _T_6391; // @[Mux.scala 27:72]
  wire [21:0] _T_6392 = _T_4974 ? _T_2141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6647 = _T_6646 | _T_6392; // @[Mux.scala 27:72]
  wire [21:0] _T_6393 = _T_4976 ? _T_2145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6648 = _T_6647 | _T_6393; // @[Mux.scala 27:72]
  wire [21:0] _T_6394 = _T_4978 ? _T_2149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6649 = _T_6648 | _T_6394; // @[Mux.scala 27:72]
  wire [21:0] _T_6395 = _T_4980 ? _T_2153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6650 = _T_6649 | _T_6395; // @[Mux.scala 27:72]
  wire [21:0] _T_6396 = _T_4982 ? _T_2157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6651 = _T_6650 | _T_6396; // @[Mux.scala 27:72]
  wire [21:0] _T_6397 = _T_4984 ? _T_2161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6652 = _T_6651 | _T_6397; // @[Mux.scala 27:72]
  wire [21:0] _T_6398 = _T_4986 ? _T_2165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6653 = _T_6652 | _T_6398; // @[Mux.scala 27:72]
  wire [21:0] _T_6399 = _T_4988 ? _T_2169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6654 = _T_6653 | _T_6399; // @[Mux.scala 27:72]
  wire [21:0] _T_6400 = _T_4990 ? _T_2173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6655 = _T_6654 | _T_6400; // @[Mux.scala 27:72]
  wire [21:0] _T_6401 = _T_4992 ? _T_2177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6656 = _T_6655 | _T_6401; // @[Mux.scala 27:72]
  wire [21:0] _T_6402 = _T_4994 ? _T_2181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6657 = _T_6656 | _T_6402; // @[Mux.scala 27:72]
  wire [21:0] _T_6403 = _T_4996 ? _T_2185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6658 = _T_6657 | _T_6403; // @[Mux.scala 27:72]
  wire [21:0] _T_6404 = _T_4998 ? _T_2189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6659 = _T_6658 | _T_6404; // @[Mux.scala 27:72]
  wire [21:0] _T_6405 = _T_5000 ? _T_2193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6660 = _T_6659 | _T_6405; // @[Mux.scala 27:72]
  wire [21:0] _T_6406 = _T_5002 ? _T_2197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6661 = _T_6660 | _T_6406; // @[Mux.scala 27:72]
  wire [21:0] _T_6407 = _T_5004 ? _T_2201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6662 = _T_6661 | _T_6407; // @[Mux.scala 27:72]
  wire [21:0] _T_6408 = _T_5006 ? _T_2205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6663 = _T_6662 | _T_6408; // @[Mux.scala 27:72]
  wire [21:0] _T_6409 = _T_5008 ? _T_2209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6664 = _T_6663 | _T_6409; // @[Mux.scala 27:72]
  wire [21:0] _T_6410 = _T_5010 ? _T_2213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6665 = _T_6664 | _T_6410; // @[Mux.scala 27:72]
  wire [21:0] _T_6411 = _T_5012 ? _T_2217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6666 = _T_6665 | _T_6411; // @[Mux.scala 27:72]
  wire [21:0] _T_6412 = _T_5014 ? _T_2221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6667 = _T_6666 | _T_6412; // @[Mux.scala 27:72]
  wire [21:0] _T_6413 = _T_5016 ? _T_2225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6668 = _T_6667 | _T_6413; // @[Mux.scala 27:72]
  wire [21:0] _T_6414 = _T_5018 ? _T_2229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6669 = _T_6668 | _T_6414; // @[Mux.scala 27:72]
  wire [21:0] _T_6415 = _T_5020 ? _T_2233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6670 = _T_6669 | _T_6415; // @[Mux.scala 27:72]
  wire [21:0] _T_6416 = _T_5022 ? _T_2237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6671 = _T_6670 | _T_6416; // @[Mux.scala 27:72]
  wire [21:0] _T_6417 = _T_5024 ? _T_2241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6672 = _T_6671 | _T_6417; // @[Mux.scala 27:72]
  wire [21:0] _T_6418 = _T_5026 ? _T_2245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6673 = _T_6672 | _T_6418; // @[Mux.scala 27:72]
  wire [21:0] _T_6419 = _T_5028 ? _T_2249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6674 = _T_6673 | _T_6419; // @[Mux.scala 27:72]
  wire [21:0] _T_6420 = _T_5030 ? _T_2253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6675 = _T_6674 | _T_6420; // @[Mux.scala 27:72]
  wire [21:0] _T_6421 = _T_5032 ? _T_2257 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6676 = _T_6675 | _T_6421; // @[Mux.scala 27:72]
  wire [21:0] _T_6422 = _T_5034 ? _T_2261 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6677 = _T_6676 | _T_6422; // @[Mux.scala 27:72]
  wire [21:0] _T_6423 = _T_5036 ? _T_2265 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6678 = _T_6677 | _T_6423; // @[Mux.scala 27:72]
  wire [21:0] _T_6424 = _T_5038 ? _T_2269 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6679 = _T_6678 | _T_6424; // @[Mux.scala 27:72]
  wire [21:0] _T_6425 = _T_5040 ? _T_2273 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6680 = _T_6679 | _T_6425; // @[Mux.scala 27:72]
  wire [21:0] _T_6426 = _T_5042 ? _T_2277 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6681 = _T_6680 | _T_6426; // @[Mux.scala 27:72]
  wire [21:0] _T_6427 = _T_5044 ? _T_2281 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6682 = _T_6681 | _T_6427; // @[Mux.scala 27:72]
  wire [21:0] _T_6428 = _T_5046 ? _T_2285 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6683 = _T_6682 | _T_6428; // @[Mux.scala 27:72]
  wire [21:0] _T_6429 = _T_5048 ? _T_2289 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6684 = _T_6683 | _T_6429; // @[Mux.scala 27:72]
  wire [21:0] _T_6430 = _T_5050 ? _T_2293 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6685 = _T_6684 | _T_6430; // @[Mux.scala 27:72]
  wire [21:0] _T_6431 = _T_5052 ? _T_2297 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6686 = _T_6685 | _T_6431; // @[Mux.scala 27:72]
  wire [21:0] _T_6432 = _T_5054 ? _T_2301 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6687 = _T_6686 | _T_6432; // @[Mux.scala 27:72]
  wire [21:0] _T_6433 = _T_5056 ? _T_2305 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6688 = _T_6687 | _T_6433; // @[Mux.scala 27:72]
  wire [21:0] _T_6434 = _T_5058 ? _T_2309 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6689 = _T_6688 | _T_6434; // @[Mux.scala 27:72]
  wire [21:0] _T_6435 = _T_5060 ? _T_2313 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6690 = _T_6689 | _T_6435; // @[Mux.scala 27:72]
  wire [21:0] _T_6436 = _T_5062 ? _T_2317 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6691 = _T_6690 | _T_6436; // @[Mux.scala 27:72]
  wire [21:0] _T_6437 = _T_5064 ? _T_2321 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6692 = _T_6691 | _T_6437; // @[Mux.scala 27:72]
  wire [21:0] _T_6438 = _T_5066 ? _T_2325 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6693 = _T_6692 | _T_6438; // @[Mux.scala 27:72]
  wire [21:0] _T_6439 = _T_5068 ? _T_2329 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6694 = _T_6693 | _T_6439; // @[Mux.scala 27:72]
  wire [21:0] _T_6440 = _T_5070 ? _T_2333 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6695 = _T_6694 | _T_6440; // @[Mux.scala 27:72]
  wire [21:0] _T_6441 = _T_5072 ? _T_2337 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6696 = _T_6695 | _T_6441; // @[Mux.scala 27:72]
  wire [21:0] _T_6442 = _T_5074 ? _T_2341 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6697 = _T_6696 | _T_6442; // @[Mux.scala 27:72]
  wire [21:0] _T_6443 = _T_5076 ? _T_2345 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6698 = _T_6697 | _T_6443; // @[Mux.scala 27:72]
  wire [21:0] _T_6444 = _T_5078 ? _T_2349 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6699 = _T_6698 | _T_6444; // @[Mux.scala 27:72]
  wire [21:0] _T_6445 = _T_5080 ? _T_2353 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6700 = _T_6699 | _T_6445; // @[Mux.scala 27:72]
  wire [21:0] _T_6446 = _T_5082 ? _T_2357 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6701 = _T_6700 | _T_6446; // @[Mux.scala 27:72]
  wire [21:0] _T_6447 = _T_5084 ? _T_2361 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6702 = _T_6701 | _T_6447; // @[Mux.scala 27:72]
  wire [21:0] _T_6448 = _T_5086 ? _T_2365 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6703 = _T_6702 | _T_6448; // @[Mux.scala 27:72]
  wire [21:0] _T_6449 = _T_5088 ? _T_2369 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6704 = _T_6703 | _T_6449; // @[Mux.scala 27:72]
  wire [21:0] _T_6450 = _T_5090 ? _T_2373 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6705 = _T_6704 | _T_6450; // @[Mux.scala 27:72]
  wire [21:0] _T_6451 = _T_5092 ? _T_2377 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6706 = _T_6705 | _T_6451; // @[Mux.scala 27:72]
  wire [21:0] _T_6452 = _T_5094 ? _T_2381 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6707 = _T_6706 | _T_6452; // @[Mux.scala 27:72]
  wire [21:0] _T_6453 = _T_5096 ? _T_2385 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6708 = _T_6707 | _T_6453; // @[Mux.scala 27:72]
  wire [21:0] _T_6454 = _T_5098 ? _T_2389 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6709 = _T_6708 | _T_6454; // @[Mux.scala 27:72]
  wire [21:0] _T_6455 = _T_5100 ? _T_2393 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6710 = _T_6709 | _T_6455; // @[Mux.scala 27:72]
  wire [21:0] _T_6456 = _T_5102 ? _T_2397 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6711 = _T_6710 | _T_6456; // @[Mux.scala 27:72]
  wire [21:0] _T_6457 = _T_5104 ? _T_2401 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6712 = _T_6711 | _T_6457; // @[Mux.scala 27:72]
  wire [21:0] _T_6458 = _T_5106 ? _T_2405 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6713 = _T_6712 | _T_6458; // @[Mux.scala 27:72]
  wire [21:0] _T_6459 = _T_5108 ? _T_2409 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6714 = _T_6713 | _T_6459; // @[Mux.scala 27:72]
  wire [21:0] _T_6460 = _T_5110 ? _T_2413 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6715 = _T_6714 | _T_6460; // @[Mux.scala 27:72]
  wire [21:0] _T_6461 = _T_5112 ? _T_2417 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6716 = _T_6715 | _T_6461; // @[Mux.scala 27:72]
  wire [21:0] _T_6462 = _T_5114 ? _T_2421 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6717 = _T_6716 | _T_6462; // @[Mux.scala 27:72]
  wire [21:0] _T_6463 = _T_5116 ? _T_2425 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6718 = _T_6717 | _T_6463; // @[Mux.scala 27:72]
  wire [21:0] _T_6464 = _T_5118 ? _T_2429 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6719 = _T_6718 | _T_6464; // @[Mux.scala 27:72]
  wire [21:0] _T_6465 = _T_5120 ? _T_2433 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6720 = _T_6719 | _T_6465; // @[Mux.scala 27:72]
  wire [21:0] _T_6466 = _T_5122 ? _T_2437 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6721 = _T_6720 | _T_6466; // @[Mux.scala 27:72]
  wire [21:0] _T_6467 = _T_5124 ? _T_2441 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6722 = _T_6721 | _T_6467; // @[Mux.scala 27:72]
  wire [21:0] _T_6468 = _T_5126 ? _T_2445 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6723 = _T_6722 | _T_6468; // @[Mux.scala 27:72]
  wire [21:0] _T_6469 = _T_5128 ? _T_2449 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6724 = _T_6723 | _T_6469; // @[Mux.scala 27:72]
  wire [21:0] _T_6470 = _T_5130 ? _T_2453 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6725 = _T_6724 | _T_6470; // @[Mux.scala 27:72]
  wire [21:0] _T_6471 = _T_5132 ? _T_2457 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6726 = _T_6725 | _T_6471; // @[Mux.scala 27:72]
  wire [21:0] _T_6472 = _T_5134 ? _T_2461 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6727 = _T_6726 | _T_6472; // @[Mux.scala 27:72]
  wire [21:0] _T_6473 = _T_5136 ? _T_2465 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6728 = _T_6727 | _T_6473; // @[Mux.scala 27:72]
  wire [21:0] _T_6474 = _T_5138 ? _T_2469 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6729 = _T_6728 | _T_6474; // @[Mux.scala 27:72]
  wire [21:0] _T_6475 = _T_5140 ? _T_2473 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6730 = _T_6729 | _T_6475; // @[Mux.scala 27:72]
  wire [21:0] _T_6476 = _T_5142 ? _T_2477 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6731 = _T_6730 | _T_6476; // @[Mux.scala 27:72]
  wire [21:0] _T_6477 = _T_5144 ? _T_2481 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6732 = _T_6731 | _T_6477; // @[Mux.scala 27:72]
  wire [21:0] _T_6478 = _T_5146 ? _T_2485 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6733 = _T_6732 | _T_6478; // @[Mux.scala 27:72]
  wire [21:0] _T_6479 = _T_5148 ? _T_2489 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6734 = _T_6733 | _T_6479; // @[Mux.scala 27:72]
  wire [21:0] _T_6480 = _T_5150 ? _T_2493 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6735 = _T_6734 | _T_6480; // @[Mux.scala 27:72]
  wire [21:0] _T_6481 = _T_5152 ? _T_2497 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6736 = _T_6735 | _T_6481; // @[Mux.scala 27:72]
  wire [21:0] _T_6482 = _T_5154 ? _T_2501 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6737 = _T_6736 | _T_6482; // @[Mux.scala 27:72]
  wire [21:0] _T_6483 = _T_5156 ? _T_2505 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6738 = _T_6737 | _T_6483; // @[Mux.scala 27:72]
  wire [21:0] _T_6484 = _T_5158 ? _T_2509 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6739 = _T_6738 | _T_6484; // @[Mux.scala 27:72]
  wire [21:0] _T_6485 = _T_5160 ? _T_2513 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6740 = _T_6739 | _T_6485; // @[Mux.scala 27:72]
  wire [21:0] _T_6486 = _T_5162 ? _T_2517 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6741 = _T_6740 | _T_6486; // @[Mux.scala 27:72]
  wire [21:0] _T_6487 = _T_5164 ? _T_2521 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6742 = _T_6741 | _T_6487; // @[Mux.scala 27:72]
  wire [21:0] _T_6488 = _T_5166 ? _T_2525 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6743 = _T_6742 | _T_6488; // @[Mux.scala 27:72]
  wire [21:0] _T_6489 = _T_5168 ? _T_2529 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6744 = _T_6743 | _T_6489; // @[Mux.scala 27:72]
  wire [21:0] _T_6490 = _T_5170 ? _T_2533 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6745 = _T_6744 | _T_6490; // @[Mux.scala 27:72]
  wire [21:0] _T_6491 = _T_5172 ? _T_2537 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6746 = _T_6745 | _T_6491; // @[Mux.scala 27:72]
  wire [21:0] _T_6492 = _T_5174 ? _T_2541 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6747 = _T_6746 | _T_6492; // @[Mux.scala 27:72]
  wire [21:0] _T_6493 = _T_5176 ? _T_2545 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6748 = _T_6747 | _T_6493; // @[Mux.scala 27:72]
  wire [21:0] _T_6494 = _T_5178 ? _T_2549 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6749 = _T_6748 | _T_6494; // @[Mux.scala 27:72]
  wire [21:0] _T_6495 = _T_5180 ? _T_2553 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6750 = _T_6749 | _T_6495; // @[Mux.scala 27:72]
  wire [21:0] _T_6496 = _T_5182 ? _T_2557 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6751 = _T_6750 | _T_6496; // @[Mux.scala 27:72]
  wire [21:0] _T_6497 = _T_5184 ? _T_2561 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6752 = _T_6751 | _T_6497; // @[Mux.scala 27:72]
  wire [21:0] _T_6498 = _T_5186 ? _T_2565 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6753 = _T_6752 | _T_6498; // @[Mux.scala 27:72]
  wire [21:0] _T_6499 = _T_5188 ? _T_2569 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6754 = _T_6753 | _T_6499; // @[Mux.scala 27:72]
  wire [21:0] _T_6500 = _T_5190 ? _T_2573 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6755 = _T_6754 | _T_6500; // @[Mux.scala 27:72]
  wire [21:0] _T_6501 = _T_5192 ? _T_2577 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6756 = _T_6755 | _T_6501; // @[Mux.scala 27:72]
  wire [21:0] _T_6502 = _T_5194 ? _T_2581 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6757 = _T_6756 | _T_6502; // @[Mux.scala 27:72]
  wire [21:0] _T_6503 = _T_5196 ? _T_2585 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6758 = _T_6757 | _T_6503; // @[Mux.scala 27:72]
  wire [21:0] _T_6504 = _T_5198 ? _T_2589 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6759 = _T_6758 | _T_6504; // @[Mux.scala 27:72]
  wire [21:0] _T_6505 = _T_5200 ? _T_2593 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6760 = _T_6759 | _T_6505; // @[Mux.scala 27:72]
  wire [21:0] _T_6506 = _T_5202 ? _T_2597 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6761 = _T_6760 | _T_6506; // @[Mux.scala 27:72]
  wire [21:0] _T_6507 = _T_5204 ? _T_2601 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6762 = _T_6761 | _T_6507; // @[Mux.scala 27:72]
  wire [21:0] _T_6508 = _T_5206 ? _T_2605 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6763 = _T_6762 | _T_6508; // @[Mux.scala 27:72]
  wire [21:0] _T_6509 = _T_5208 ? _T_2609 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6764 = _T_6763 | _T_6509; // @[Mux.scala 27:72]
  wire [21:0] _T_6510 = _T_5210 ? _T_2613 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6765 = _T_6764 | _T_6510; // @[Mux.scala 27:72]
  wire [21:0] _T_6511 = _T_5212 ? _T_2617 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6766 = _T_6765 | _T_6511; // @[Mux.scala 27:72]
  wire [21:0] _T_6512 = _T_5214 ? _T_2621 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6767 = _T_6766 | _T_6512; // @[Mux.scala 27:72]
  wire [21:0] _T_6513 = _T_5216 ? _T_2625 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6768 = _T_6767 | _T_6513; // @[Mux.scala 27:72]
  wire [21:0] _T_6514 = _T_5218 ? _T_2629 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6769 = _T_6768 | _T_6514; // @[Mux.scala 27:72]
  wire [21:0] _T_6515 = _T_5220 ? _T_2633 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6770 = _T_6769 | _T_6515; // @[Mux.scala 27:72]
  wire [21:0] _T_6516 = _T_5222 ? _T_2637 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6771 = _T_6770 | _T_6516; // @[Mux.scala 27:72]
  wire [21:0] _T_6517 = _T_5224 ? _T_2641 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6772 = _T_6771 | _T_6517; // @[Mux.scala 27:72]
  wire [21:0] _T_6518 = _T_5226 ? _T_2645 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6773 = _T_6772 | _T_6518; // @[Mux.scala 27:72]
  wire [21:0] _T_6519 = _T_5228 ? _T_2649 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6774 = _T_6773 | _T_6519; // @[Mux.scala 27:72]
  wire [21:0] _T_6520 = _T_5230 ? _T_2653 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6775 = _T_6774 | _T_6520; // @[Mux.scala 27:72]
  wire [21:0] _T_6521 = _T_5232 ? _T_2657 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6776 = _T_6775 | _T_6521; // @[Mux.scala 27:72]
  wire [21:0] _T_6522 = _T_5234 ? _T_2661 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6777 = _T_6776 | _T_6522; // @[Mux.scala 27:72]
  wire [21:0] _T_6523 = _T_5236 ? _T_2665 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6778 = _T_6777 | _T_6523; // @[Mux.scala 27:72]
  wire [21:0] _T_6524 = _T_5238 ? _T_2669 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6779 = _T_6778 | _T_6524; // @[Mux.scala 27:72]
  wire [21:0] _T_6525 = _T_5240 ? _T_2673 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6780 = _T_6779 | _T_6525; // @[Mux.scala 27:72]
  wire [21:0] _T_6526 = _T_5242 ? _T_2677 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6781 = _T_6780 | _T_6526; // @[Mux.scala 27:72]
  wire [21:0] _T_6527 = _T_5244 ? _T_2681 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6782 = _T_6781 | _T_6527; // @[Mux.scala 27:72]
  wire [21:0] _T_6528 = _T_5246 ? _T_2685 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6783 = _T_6782 | _T_6528; // @[Mux.scala 27:72]
  wire [21:0] _T_6529 = _T_5248 ? _T_2689 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6784 = _T_6783 | _T_6529; // @[Mux.scala 27:72]
  wire [21:0] _T_6785 = _T_6784; // @[Mux.scala 27:72 Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_p1_f = _T_6784; // @[ifu_bp_ctl.scala 444:31]
  wire  _T_80 = _T_6785[21:17] == _T_37; // @[ifu_bp_ctl.scala 155:107]
  wire  _T_81 = _T_6785[0] & _T_80; // @[ifu_bp_ctl.scala 155:61]
  wire  _T_84 = _T_81 & _T_73; // @[ifu_bp_ctl.scala 155:130]
  wire  _T_85 = _T_84 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 156:57]
  wire  _T_87 = _T_85 & _T; // @[ifu_bp_ctl.scala 156:78]
  wire  _T_120 = _T_6785[3] ^ _T_6785[4]; // @[ifu_bp_ctl.scala 168:99]
  wire  _T_121 = _T_87 & _T_120; // @[ifu_bp_ctl.scala 168:62]
  wire  _T_125 = ~_T_120; // @[ifu_bp_ctl.scala 169:27]
  wire  _T_126 = _T_87 & _T_125; // @[ifu_bp_ctl.scala 169:25]
  wire [1:0] _T_127 = {_T_121,_T_126}; // @[Cat.scala 29:58]
  wire [21:0] _T_151 = _T_127[0] ? _T_6785 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_152 = _T_150 | _T_151; // @[Mux.scala 27:72]
  wire [21:0] _T_165 = io_ifc_fetch_addr_f[0] ? _T_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank1_rd_data_f = _T_164 | _T_165; // @[Mux.scala 27:72]
  wire  _T_262 = btb_vbank1_rd_data_f[2] | btb_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 280:59]
  wire [21:0] _T_134 = _T_97[0] ? _T_3713 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_135 = _T_107[0] ? _T_4737 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_136 = _T_134 | _T_135; // @[Mux.scala 27:72]
  wire [21:0] _T_157 = _T_162 ? _T_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_158 = io_ifc_fetch_addr_f[0] ? _T_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank0_rd_data_f = _T_157 | _T_158; // @[Mux.scala 27:72]
  wire  _T_265 = btb_vbank0_rd_data_f[2] | btb_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 281:59]
  wire [1:0] bht_force_taken_f = {_T_262,_T_265}; // @[Cat.scala 29:58]
  wire [9:0] _T_608 = {btb_rd_addr_f,2'h0}; // @[Cat.scala 29:58]
  reg [7:0] fghr; // @[Reg.scala 27:20]
  wire [7:0] bht_rd_addr_f = _T_608[9:2] ^ fghr; // @[lib.scala 56:35]
  wire  _T_22498 = bht_rd_addr_f == 8'h0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_0; // @[Reg.scala 27:20]
  wire [1:0] _T_23010 = _T_22498 ? bht_bank_rd_data_out_1_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_22500 = bht_rd_addr_f == 8'h1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_1; // @[Reg.scala 27:20]
  wire [1:0] _T_23011 = _T_22500 ? bht_bank_rd_data_out_1_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23266 = _T_23010 | _T_23011; // @[Mux.scala 27:72]
  wire  _T_22502 = bht_rd_addr_f == 8'h2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_2; // @[Reg.scala 27:20]
  wire [1:0] _T_23012 = _T_22502 ? bht_bank_rd_data_out_1_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23267 = _T_23266 | _T_23012; // @[Mux.scala 27:72]
  wire  _T_22504 = bht_rd_addr_f == 8'h3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_3; // @[Reg.scala 27:20]
  wire [1:0] _T_23013 = _T_22504 ? bht_bank_rd_data_out_1_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23268 = _T_23267 | _T_23013; // @[Mux.scala 27:72]
  wire  _T_22506 = bht_rd_addr_f == 8'h4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_4; // @[Reg.scala 27:20]
  wire [1:0] _T_23014 = _T_22506 ? bht_bank_rd_data_out_1_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23269 = _T_23268 | _T_23014; // @[Mux.scala 27:72]
  wire  _T_22508 = bht_rd_addr_f == 8'h5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_5; // @[Reg.scala 27:20]
  wire [1:0] _T_23015 = _T_22508 ? bht_bank_rd_data_out_1_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23270 = _T_23269 | _T_23015; // @[Mux.scala 27:72]
  wire  _T_22510 = bht_rd_addr_f == 8'h6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_6; // @[Reg.scala 27:20]
  wire [1:0] _T_23016 = _T_22510 ? bht_bank_rd_data_out_1_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23271 = _T_23270 | _T_23016; // @[Mux.scala 27:72]
  wire  _T_22512 = bht_rd_addr_f == 8'h7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_7; // @[Reg.scala 27:20]
  wire [1:0] _T_23017 = _T_22512 ? bht_bank_rd_data_out_1_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23272 = _T_23271 | _T_23017; // @[Mux.scala 27:72]
  wire  _T_22514 = bht_rd_addr_f == 8'h8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_8; // @[Reg.scala 27:20]
  wire [1:0] _T_23018 = _T_22514 ? bht_bank_rd_data_out_1_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23273 = _T_23272 | _T_23018; // @[Mux.scala 27:72]
  wire  _T_22516 = bht_rd_addr_f == 8'h9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_9; // @[Reg.scala 27:20]
  wire [1:0] _T_23019 = _T_22516 ? bht_bank_rd_data_out_1_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23274 = _T_23273 | _T_23019; // @[Mux.scala 27:72]
  wire  _T_22518 = bht_rd_addr_f == 8'ha; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_10; // @[Reg.scala 27:20]
  wire [1:0] _T_23020 = _T_22518 ? bht_bank_rd_data_out_1_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23275 = _T_23274 | _T_23020; // @[Mux.scala 27:72]
  wire  _T_22520 = bht_rd_addr_f == 8'hb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_11; // @[Reg.scala 27:20]
  wire [1:0] _T_23021 = _T_22520 ? bht_bank_rd_data_out_1_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23276 = _T_23275 | _T_23021; // @[Mux.scala 27:72]
  wire  _T_22522 = bht_rd_addr_f == 8'hc; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_12; // @[Reg.scala 27:20]
  wire [1:0] _T_23022 = _T_22522 ? bht_bank_rd_data_out_1_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23277 = _T_23276 | _T_23022; // @[Mux.scala 27:72]
  wire  _T_22524 = bht_rd_addr_f == 8'hd; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_13; // @[Reg.scala 27:20]
  wire [1:0] _T_23023 = _T_22524 ? bht_bank_rd_data_out_1_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23278 = _T_23277 | _T_23023; // @[Mux.scala 27:72]
  wire  _T_22526 = bht_rd_addr_f == 8'he; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_14; // @[Reg.scala 27:20]
  wire [1:0] _T_23024 = _T_22526 ? bht_bank_rd_data_out_1_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23279 = _T_23278 | _T_23024; // @[Mux.scala 27:72]
  wire  _T_22528 = bht_rd_addr_f == 8'hf; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_15; // @[Reg.scala 27:20]
  wire [1:0] _T_23025 = _T_22528 ? bht_bank_rd_data_out_1_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23280 = _T_23279 | _T_23025; // @[Mux.scala 27:72]
  wire  _T_22530 = bht_rd_addr_f == 8'h10; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_16; // @[Reg.scala 27:20]
  wire [1:0] _T_23026 = _T_22530 ? bht_bank_rd_data_out_1_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23281 = _T_23280 | _T_23026; // @[Mux.scala 27:72]
  wire  _T_22532 = bht_rd_addr_f == 8'h11; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_17; // @[Reg.scala 27:20]
  wire [1:0] _T_23027 = _T_22532 ? bht_bank_rd_data_out_1_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23282 = _T_23281 | _T_23027; // @[Mux.scala 27:72]
  wire  _T_22534 = bht_rd_addr_f == 8'h12; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_18; // @[Reg.scala 27:20]
  wire [1:0] _T_23028 = _T_22534 ? bht_bank_rd_data_out_1_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23283 = _T_23282 | _T_23028; // @[Mux.scala 27:72]
  wire  _T_22536 = bht_rd_addr_f == 8'h13; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_19; // @[Reg.scala 27:20]
  wire [1:0] _T_23029 = _T_22536 ? bht_bank_rd_data_out_1_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23284 = _T_23283 | _T_23029; // @[Mux.scala 27:72]
  wire  _T_22538 = bht_rd_addr_f == 8'h14; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_20; // @[Reg.scala 27:20]
  wire [1:0] _T_23030 = _T_22538 ? bht_bank_rd_data_out_1_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23285 = _T_23284 | _T_23030; // @[Mux.scala 27:72]
  wire  _T_22540 = bht_rd_addr_f == 8'h15; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_21; // @[Reg.scala 27:20]
  wire [1:0] _T_23031 = _T_22540 ? bht_bank_rd_data_out_1_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23286 = _T_23285 | _T_23031; // @[Mux.scala 27:72]
  wire  _T_22542 = bht_rd_addr_f == 8'h16; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_22; // @[Reg.scala 27:20]
  wire [1:0] _T_23032 = _T_22542 ? bht_bank_rd_data_out_1_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23287 = _T_23286 | _T_23032; // @[Mux.scala 27:72]
  wire  _T_22544 = bht_rd_addr_f == 8'h17; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_23; // @[Reg.scala 27:20]
  wire [1:0] _T_23033 = _T_22544 ? bht_bank_rd_data_out_1_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23288 = _T_23287 | _T_23033; // @[Mux.scala 27:72]
  wire  _T_22546 = bht_rd_addr_f == 8'h18; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_24; // @[Reg.scala 27:20]
  wire [1:0] _T_23034 = _T_22546 ? bht_bank_rd_data_out_1_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23289 = _T_23288 | _T_23034; // @[Mux.scala 27:72]
  wire  _T_22548 = bht_rd_addr_f == 8'h19; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_25; // @[Reg.scala 27:20]
  wire [1:0] _T_23035 = _T_22548 ? bht_bank_rd_data_out_1_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23290 = _T_23289 | _T_23035; // @[Mux.scala 27:72]
  wire  _T_22550 = bht_rd_addr_f == 8'h1a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_26; // @[Reg.scala 27:20]
  wire [1:0] _T_23036 = _T_22550 ? bht_bank_rd_data_out_1_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23291 = _T_23290 | _T_23036; // @[Mux.scala 27:72]
  wire  _T_22552 = bht_rd_addr_f == 8'h1b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_27; // @[Reg.scala 27:20]
  wire [1:0] _T_23037 = _T_22552 ? bht_bank_rd_data_out_1_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23292 = _T_23291 | _T_23037; // @[Mux.scala 27:72]
  wire  _T_22554 = bht_rd_addr_f == 8'h1c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_28; // @[Reg.scala 27:20]
  wire [1:0] _T_23038 = _T_22554 ? bht_bank_rd_data_out_1_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23293 = _T_23292 | _T_23038; // @[Mux.scala 27:72]
  wire  _T_22556 = bht_rd_addr_f == 8'h1d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_29; // @[Reg.scala 27:20]
  wire [1:0] _T_23039 = _T_22556 ? bht_bank_rd_data_out_1_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23294 = _T_23293 | _T_23039; // @[Mux.scala 27:72]
  wire  _T_22558 = bht_rd_addr_f == 8'h1e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_30; // @[Reg.scala 27:20]
  wire [1:0] _T_23040 = _T_22558 ? bht_bank_rd_data_out_1_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23295 = _T_23294 | _T_23040; // @[Mux.scala 27:72]
  wire  _T_22560 = bht_rd_addr_f == 8'h1f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_31; // @[Reg.scala 27:20]
  wire [1:0] _T_23041 = _T_22560 ? bht_bank_rd_data_out_1_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23296 = _T_23295 | _T_23041; // @[Mux.scala 27:72]
  wire  _T_22562 = bht_rd_addr_f == 8'h20; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_32; // @[Reg.scala 27:20]
  wire [1:0] _T_23042 = _T_22562 ? bht_bank_rd_data_out_1_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23297 = _T_23296 | _T_23042; // @[Mux.scala 27:72]
  wire  _T_22564 = bht_rd_addr_f == 8'h21; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_33; // @[Reg.scala 27:20]
  wire [1:0] _T_23043 = _T_22564 ? bht_bank_rd_data_out_1_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23298 = _T_23297 | _T_23043; // @[Mux.scala 27:72]
  wire  _T_22566 = bht_rd_addr_f == 8'h22; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_34; // @[Reg.scala 27:20]
  wire [1:0] _T_23044 = _T_22566 ? bht_bank_rd_data_out_1_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23299 = _T_23298 | _T_23044; // @[Mux.scala 27:72]
  wire  _T_22568 = bht_rd_addr_f == 8'h23; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_35; // @[Reg.scala 27:20]
  wire [1:0] _T_23045 = _T_22568 ? bht_bank_rd_data_out_1_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23300 = _T_23299 | _T_23045; // @[Mux.scala 27:72]
  wire  _T_22570 = bht_rd_addr_f == 8'h24; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_36; // @[Reg.scala 27:20]
  wire [1:0] _T_23046 = _T_22570 ? bht_bank_rd_data_out_1_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23301 = _T_23300 | _T_23046; // @[Mux.scala 27:72]
  wire  _T_22572 = bht_rd_addr_f == 8'h25; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_37; // @[Reg.scala 27:20]
  wire [1:0] _T_23047 = _T_22572 ? bht_bank_rd_data_out_1_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23302 = _T_23301 | _T_23047; // @[Mux.scala 27:72]
  wire  _T_22574 = bht_rd_addr_f == 8'h26; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_38; // @[Reg.scala 27:20]
  wire [1:0] _T_23048 = _T_22574 ? bht_bank_rd_data_out_1_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23303 = _T_23302 | _T_23048; // @[Mux.scala 27:72]
  wire  _T_22576 = bht_rd_addr_f == 8'h27; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_39; // @[Reg.scala 27:20]
  wire [1:0] _T_23049 = _T_22576 ? bht_bank_rd_data_out_1_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23304 = _T_23303 | _T_23049; // @[Mux.scala 27:72]
  wire  _T_22578 = bht_rd_addr_f == 8'h28; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_40; // @[Reg.scala 27:20]
  wire [1:0] _T_23050 = _T_22578 ? bht_bank_rd_data_out_1_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23305 = _T_23304 | _T_23050; // @[Mux.scala 27:72]
  wire  _T_22580 = bht_rd_addr_f == 8'h29; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_41; // @[Reg.scala 27:20]
  wire [1:0] _T_23051 = _T_22580 ? bht_bank_rd_data_out_1_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23306 = _T_23305 | _T_23051; // @[Mux.scala 27:72]
  wire  _T_22582 = bht_rd_addr_f == 8'h2a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_42; // @[Reg.scala 27:20]
  wire [1:0] _T_23052 = _T_22582 ? bht_bank_rd_data_out_1_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23307 = _T_23306 | _T_23052; // @[Mux.scala 27:72]
  wire  _T_22584 = bht_rd_addr_f == 8'h2b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_43; // @[Reg.scala 27:20]
  wire [1:0] _T_23053 = _T_22584 ? bht_bank_rd_data_out_1_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23308 = _T_23307 | _T_23053; // @[Mux.scala 27:72]
  wire  _T_22586 = bht_rd_addr_f == 8'h2c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_44; // @[Reg.scala 27:20]
  wire [1:0] _T_23054 = _T_22586 ? bht_bank_rd_data_out_1_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23309 = _T_23308 | _T_23054; // @[Mux.scala 27:72]
  wire  _T_22588 = bht_rd_addr_f == 8'h2d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_45; // @[Reg.scala 27:20]
  wire [1:0] _T_23055 = _T_22588 ? bht_bank_rd_data_out_1_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23310 = _T_23309 | _T_23055; // @[Mux.scala 27:72]
  wire  _T_22590 = bht_rd_addr_f == 8'h2e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_46; // @[Reg.scala 27:20]
  wire [1:0] _T_23056 = _T_22590 ? bht_bank_rd_data_out_1_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23311 = _T_23310 | _T_23056; // @[Mux.scala 27:72]
  wire  _T_22592 = bht_rd_addr_f == 8'h2f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_47; // @[Reg.scala 27:20]
  wire [1:0] _T_23057 = _T_22592 ? bht_bank_rd_data_out_1_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23312 = _T_23311 | _T_23057; // @[Mux.scala 27:72]
  wire  _T_22594 = bht_rd_addr_f == 8'h30; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_48; // @[Reg.scala 27:20]
  wire [1:0] _T_23058 = _T_22594 ? bht_bank_rd_data_out_1_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23313 = _T_23312 | _T_23058; // @[Mux.scala 27:72]
  wire  _T_22596 = bht_rd_addr_f == 8'h31; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_49; // @[Reg.scala 27:20]
  wire [1:0] _T_23059 = _T_22596 ? bht_bank_rd_data_out_1_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23314 = _T_23313 | _T_23059; // @[Mux.scala 27:72]
  wire  _T_22598 = bht_rd_addr_f == 8'h32; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_50; // @[Reg.scala 27:20]
  wire [1:0] _T_23060 = _T_22598 ? bht_bank_rd_data_out_1_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23315 = _T_23314 | _T_23060; // @[Mux.scala 27:72]
  wire  _T_22600 = bht_rd_addr_f == 8'h33; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_51; // @[Reg.scala 27:20]
  wire [1:0] _T_23061 = _T_22600 ? bht_bank_rd_data_out_1_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23316 = _T_23315 | _T_23061; // @[Mux.scala 27:72]
  wire  _T_22602 = bht_rd_addr_f == 8'h34; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_52; // @[Reg.scala 27:20]
  wire [1:0] _T_23062 = _T_22602 ? bht_bank_rd_data_out_1_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23317 = _T_23316 | _T_23062; // @[Mux.scala 27:72]
  wire  _T_22604 = bht_rd_addr_f == 8'h35; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_53; // @[Reg.scala 27:20]
  wire [1:0] _T_23063 = _T_22604 ? bht_bank_rd_data_out_1_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23318 = _T_23317 | _T_23063; // @[Mux.scala 27:72]
  wire  _T_22606 = bht_rd_addr_f == 8'h36; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_54; // @[Reg.scala 27:20]
  wire [1:0] _T_23064 = _T_22606 ? bht_bank_rd_data_out_1_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23319 = _T_23318 | _T_23064; // @[Mux.scala 27:72]
  wire  _T_22608 = bht_rd_addr_f == 8'h37; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_55; // @[Reg.scala 27:20]
  wire [1:0] _T_23065 = _T_22608 ? bht_bank_rd_data_out_1_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23320 = _T_23319 | _T_23065; // @[Mux.scala 27:72]
  wire  _T_22610 = bht_rd_addr_f == 8'h38; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_56; // @[Reg.scala 27:20]
  wire [1:0] _T_23066 = _T_22610 ? bht_bank_rd_data_out_1_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23321 = _T_23320 | _T_23066; // @[Mux.scala 27:72]
  wire  _T_22612 = bht_rd_addr_f == 8'h39; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_57; // @[Reg.scala 27:20]
  wire [1:0] _T_23067 = _T_22612 ? bht_bank_rd_data_out_1_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23322 = _T_23321 | _T_23067; // @[Mux.scala 27:72]
  wire  _T_22614 = bht_rd_addr_f == 8'h3a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_58; // @[Reg.scala 27:20]
  wire [1:0] _T_23068 = _T_22614 ? bht_bank_rd_data_out_1_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23323 = _T_23322 | _T_23068; // @[Mux.scala 27:72]
  wire  _T_22616 = bht_rd_addr_f == 8'h3b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_59; // @[Reg.scala 27:20]
  wire [1:0] _T_23069 = _T_22616 ? bht_bank_rd_data_out_1_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23324 = _T_23323 | _T_23069; // @[Mux.scala 27:72]
  wire  _T_22618 = bht_rd_addr_f == 8'h3c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_60; // @[Reg.scala 27:20]
  wire [1:0] _T_23070 = _T_22618 ? bht_bank_rd_data_out_1_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23325 = _T_23324 | _T_23070; // @[Mux.scala 27:72]
  wire  _T_22620 = bht_rd_addr_f == 8'h3d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_61; // @[Reg.scala 27:20]
  wire [1:0] _T_23071 = _T_22620 ? bht_bank_rd_data_out_1_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23326 = _T_23325 | _T_23071; // @[Mux.scala 27:72]
  wire  _T_22622 = bht_rd_addr_f == 8'h3e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_62; // @[Reg.scala 27:20]
  wire [1:0] _T_23072 = _T_22622 ? bht_bank_rd_data_out_1_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23327 = _T_23326 | _T_23072; // @[Mux.scala 27:72]
  wire  _T_22624 = bht_rd_addr_f == 8'h3f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_63; // @[Reg.scala 27:20]
  wire [1:0] _T_23073 = _T_22624 ? bht_bank_rd_data_out_1_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23328 = _T_23327 | _T_23073; // @[Mux.scala 27:72]
  wire  _T_22626 = bht_rd_addr_f == 8'h40; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_64; // @[Reg.scala 27:20]
  wire [1:0] _T_23074 = _T_22626 ? bht_bank_rd_data_out_1_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23329 = _T_23328 | _T_23074; // @[Mux.scala 27:72]
  wire  _T_22628 = bht_rd_addr_f == 8'h41; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_65; // @[Reg.scala 27:20]
  wire [1:0] _T_23075 = _T_22628 ? bht_bank_rd_data_out_1_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23330 = _T_23329 | _T_23075; // @[Mux.scala 27:72]
  wire  _T_22630 = bht_rd_addr_f == 8'h42; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_66; // @[Reg.scala 27:20]
  wire [1:0] _T_23076 = _T_22630 ? bht_bank_rd_data_out_1_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23331 = _T_23330 | _T_23076; // @[Mux.scala 27:72]
  wire  _T_22632 = bht_rd_addr_f == 8'h43; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_67; // @[Reg.scala 27:20]
  wire [1:0] _T_23077 = _T_22632 ? bht_bank_rd_data_out_1_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23332 = _T_23331 | _T_23077; // @[Mux.scala 27:72]
  wire  _T_22634 = bht_rd_addr_f == 8'h44; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_68; // @[Reg.scala 27:20]
  wire [1:0] _T_23078 = _T_22634 ? bht_bank_rd_data_out_1_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23333 = _T_23332 | _T_23078; // @[Mux.scala 27:72]
  wire  _T_22636 = bht_rd_addr_f == 8'h45; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_69; // @[Reg.scala 27:20]
  wire [1:0] _T_23079 = _T_22636 ? bht_bank_rd_data_out_1_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23334 = _T_23333 | _T_23079; // @[Mux.scala 27:72]
  wire  _T_22638 = bht_rd_addr_f == 8'h46; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_70; // @[Reg.scala 27:20]
  wire [1:0] _T_23080 = _T_22638 ? bht_bank_rd_data_out_1_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23335 = _T_23334 | _T_23080; // @[Mux.scala 27:72]
  wire  _T_22640 = bht_rd_addr_f == 8'h47; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_71; // @[Reg.scala 27:20]
  wire [1:0] _T_23081 = _T_22640 ? bht_bank_rd_data_out_1_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23336 = _T_23335 | _T_23081; // @[Mux.scala 27:72]
  wire  _T_22642 = bht_rd_addr_f == 8'h48; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_72; // @[Reg.scala 27:20]
  wire [1:0] _T_23082 = _T_22642 ? bht_bank_rd_data_out_1_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23337 = _T_23336 | _T_23082; // @[Mux.scala 27:72]
  wire  _T_22644 = bht_rd_addr_f == 8'h49; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_73; // @[Reg.scala 27:20]
  wire [1:0] _T_23083 = _T_22644 ? bht_bank_rd_data_out_1_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23338 = _T_23337 | _T_23083; // @[Mux.scala 27:72]
  wire  _T_22646 = bht_rd_addr_f == 8'h4a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_74; // @[Reg.scala 27:20]
  wire [1:0] _T_23084 = _T_22646 ? bht_bank_rd_data_out_1_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23339 = _T_23338 | _T_23084; // @[Mux.scala 27:72]
  wire  _T_22648 = bht_rd_addr_f == 8'h4b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_75; // @[Reg.scala 27:20]
  wire [1:0] _T_23085 = _T_22648 ? bht_bank_rd_data_out_1_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23340 = _T_23339 | _T_23085; // @[Mux.scala 27:72]
  wire  _T_22650 = bht_rd_addr_f == 8'h4c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_76; // @[Reg.scala 27:20]
  wire [1:0] _T_23086 = _T_22650 ? bht_bank_rd_data_out_1_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23341 = _T_23340 | _T_23086; // @[Mux.scala 27:72]
  wire  _T_22652 = bht_rd_addr_f == 8'h4d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_77; // @[Reg.scala 27:20]
  wire [1:0] _T_23087 = _T_22652 ? bht_bank_rd_data_out_1_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23342 = _T_23341 | _T_23087; // @[Mux.scala 27:72]
  wire  _T_22654 = bht_rd_addr_f == 8'h4e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_78; // @[Reg.scala 27:20]
  wire [1:0] _T_23088 = _T_22654 ? bht_bank_rd_data_out_1_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23343 = _T_23342 | _T_23088; // @[Mux.scala 27:72]
  wire  _T_22656 = bht_rd_addr_f == 8'h4f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_79; // @[Reg.scala 27:20]
  wire [1:0] _T_23089 = _T_22656 ? bht_bank_rd_data_out_1_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23344 = _T_23343 | _T_23089; // @[Mux.scala 27:72]
  wire  _T_22658 = bht_rd_addr_f == 8'h50; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_80; // @[Reg.scala 27:20]
  wire [1:0] _T_23090 = _T_22658 ? bht_bank_rd_data_out_1_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23345 = _T_23344 | _T_23090; // @[Mux.scala 27:72]
  wire  _T_22660 = bht_rd_addr_f == 8'h51; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_81; // @[Reg.scala 27:20]
  wire [1:0] _T_23091 = _T_22660 ? bht_bank_rd_data_out_1_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23346 = _T_23345 | _T_23091; // @[Mux.scala 27:72]
  wire  _T_22662 = bht_rd_addr_f == 8'h52; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_82; // @[Reg.scala 27:20]
  wire [1:0] _T_23092 = _T_22662 ? bht_bank_rd_data_out_1_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23347 = _T_23346 | _T_23092; // @[Mux.scala 27:72]
  wire  _T_22664 = bht_rd_addr_f == 8'h53; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_83; // @[Reg.scala 27:20]
  wire [1:0] _T_23093 = _T_22664 ? bht_bank_rd_data_out_1_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23348 = _T_23347 | _T_23093; // @[Mux.scala 27:72]
  wire  _T_22666 = bht_rd_addr_f == 8'h54; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_84; // @[Reg.scala 27:20]
  wire [1:0] _T_23094 = _T_22666 ? bht_bank_rd_data_out_1_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23349 = _T_23348 | _T_23094; // @[Mux.scala 27:72]
  wire  _T_22668 = bht_rd_addr_f == 8'h55; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_85; // @[Reg.scala 27:20]
  wire [1:0] _T_23095 = _T_22668 ? bht_bank_rd_data_out_1_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23350 = _T_23349 | _T_23095; // @[Mux.scala 27:72]
  wire  _T_22670 = bht_rd_addr_f == 8'h56; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_86; // @[Reg.scala 27:20]
  wire [1:0] _T_23096 = _T_22670 ? bht_bank_rd_data_out_1_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23351 = _T_23350 | _T_23096; // @[Mux.scala 27:72]
  wire  _T_22672 = bht_rd_addr_f == 8'h57; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_87; // @[Reg.scala 27:20]
  wire [1:0] _T_23097 = _T_22672 ? bht_bank_rd_data_out_1_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23352 = _T_23351 | _T_23097; // @[Mux.scala 27:72]
  wire  _T_22674 = bht_rd_addr_f == 8'h58; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_88; // @[Reg.scala 27:20]
  wire [1:0] _T_23098 = _T_22674 ? bht_bank_rd_data_out_1_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23353 = _T_23352 | _T_23098; // @[Mux.scala 27:72]
  wire  _T_22676 = bht_rd_addr_f == 8'h59; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_89; // @[Reg.scala 27:20]
  wire [1:0] _T_23099 = _T_22676 ? bht_bank_rd_data_out_1_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23354 = _T_23353 | _T_23099; // @[Mux.scala 27:72]
  wire  _T_22678 = bht_rd_addr_f == 8'h5a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_90; // @[Reg.scala 27:20]
  wire [1:0] _T_23100 = _T_22678 ? bht_bank_rd_data_out_1_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23355 = _T_23354 | _T_23100; // @[Mux.scala 27:72]
  wire  _T_22680 = bht_rd_addr_f == 8'h5b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_91; // @[Reg.scala 27:20]
  wire [1:0] _T_23101 = _T_22680 ? bht_bank_rd_data_out_1_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23356 = _T_23355 | _T_23101; // @[Mux.scala 27:72]
  wire  _T_22682 = bht_rd_addr_f == 8'h5c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_92; // @[Reg.scala 27:20]
  wire [1:0] _T_23102 = _T_22682 ? bht_bank_rd_data_out_1_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23357 = _T_23356 | _T_23102; // @[Mux.scala 27:72]
  wire  _T_22684 = bht_rd_addr_f == 8'h5d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_93; // @[Reg.scala 27:20]
  wire [1:0] _T_23103 = _T_22684 ? bht_bank_rd_data_out_1_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23358 = _T_23357 | _T_23103; // @[Mux.scala 27:72]
  wire  _T_22686 = bht_rd_addr_f == 8'h5e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_94; // @[Reg.scala 27:20]
  wire [1:0] _T_23104 = _T_22686 ? bht_bank_rd_data_out_1_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23359 = _T_23358 | _T_23104; // @[Mux.scala 27:72]
  wire  _T_22688 = bht_rd_addr_f == 8'h5f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_95; // @[Reg.scala 27:20]
  wire [1:0] _T_23105 = _T_22688 ? bht_bank_rd_data_out_1_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23360 = _T_23359 | _T_23105; // @[Mux.scala 27:72]
  wire  _T_22690 = bht_rd_addr_f == 8'h60; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_96; // @[Reg.scala 27:20]
  wire [1:0] _T_23106 = _T_22690 ? bht_bank_rd_data_out_1_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23361 = _T_23360 | _T_23106; // @[Mux.scala 27:72]
  wire  _T_22692 = bht_rd_addr_f == 8'h61; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_97; // @[Reg.scala 27:20]
  wire [1:0] _T_23107 = _T_22692 ? bht_bank_rd_data_out_1_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23362 = _T_23361 | _T_23107; // @[Mux.scala 27:72]
  wire  _T_22694 = bht_rd_addr_f == 8'h62; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_98; // @[Reg.scala 27:20]
  wire [1:0] _T_23108 = _T_22694 ? bht_bank_rd_data_out_1_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23363 = _T_23362 | _T_23108; // @[Mux.scala 27:72]
  wire  _T_22696 = bht_rd_addr_f == 8'h63; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_99; // @[Reg.scala 27:20]
  wire [1:0] _T_23109 = _T_22696 ? bht_bank_rd_data_out_1_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23364 = _T_23363 | _T_23109; // @[Mux.scala 27:72]
  wire  _T_22698 = bht_rd_addr_f == 8'h64; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_100; // @[Reg.scala 27:20]
  wire [1:0] _T_23110 = _T_22698 ? bht_bank_rd_data_out_1_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23365 = _T_23364 | _T_23110; // @[Mux.scala 27:72]
  wire  _T_22700 = bht_rd_addr_f == 8'h65; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_101; // @[Reg.scala 27:20]
  wire [1:0] _T_23111 = _T_22700 ? bht_bank_rd_data_out_1_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23366 = _T_23365 | _T_23111; // @[Mux.scala 27:72]
  wire  _T_22702 = bht_rd_addr_f == 8'h66; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_102; // @[Reg.scala 27:20]
  wire [1:0] _T_23112 = _T_22702 ? bht_bank_rd_data_out_1_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23367 = _T_23366 | _T_23112; // @[Mux.scala 27:72]
  wire  _T_22704 = bht_rd_addr_f == 8'h67; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_103; // @[Reg.scala 27:20]
  wire [1:0] _T_23113 = _T_22704 ? bht_bank_rd_data_out_1_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23368 = _T_23367 | _T_23113; // @[Mux.scala 27:72]
  wire  _T_22706 = bht_rd_addr_f == 8'h68; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_104; // @[Reg.scala 27:20]
  wire [1:0] _T_23114 = _T_22706 ? bht_bank_rd_data_out_1_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23369 = _T_23368 | _T_23114; // @[Mux.scala 27:72]
  wire  _T_22708 = bht_rd_addr_f == 8'h69; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_105; // @[Reg.scala 27:20]
  wire [1:0] _T_23115 = _T_22708 ? bht_bank_rd_data_out_1_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23370 = _T_23369 | _T_23115; // @[Mux.scala 27:72]
  wire  _T_22710 = bht_rd_addr_f == 8'h6a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_106; // @[Reg.scala 27:20]
  wire [1:0] _T_23116 = _T_22710 ? bht_bank_rd_data_out_1_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23371 = _T_23370 | _T_23116; // @[Mux.scala 27:72]
  wire  _T_22712 = bht_rd_addr_f == 8'h6b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_107; // @[Reg.scala 27:20]
  wire [1:0] _T_23117 = _T_22712 ? bht_bank_rd_data_out_1_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23372 = _T_23371 | _T_23117; // @[Mux.scala 27:72]
  wire  _T_22714 = bht_rd_addr_f == 8'h6c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_108; // @[Reg.scala 27:20]
  wire [1:0] _T_23118 = _T_22714 ? bht_bank_rd_data_out_1_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23373 = _T_23372 | _T_23118; // @[Mux.scala 27:72]
  wire  _T_22716 = bht_rd_addr_f == 8'h6d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_109; // @[Reg.scala 27:20]
  wire [1:0] _T_23119 = _T_22716 ? bht_bank_rd_data_out_1_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23374 = _T_23373 | _T_23119; // @[Mux.scala 27:72]
  wire  _T_22718 = bht_rd_addr_f == 8'h6e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_110; // @[Reg.scala 27:20]
  wire [1:0] _T_23120 = _T_22718 ? bht_bank_rd_data_out_1_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23375 = _T_23374 | _T_23120; // @[Mux.scala 27:72]
  wire  _T_22720 = bht_rd_addr_f == 8'h6f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_111; // @[Reg.scala 27:20]
  wire [1:0] _T_23121 = _T_22720 ? bht_bank_rd_data_out_1_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23376 = _T_23375 | _T_23121; // @[Mux.scala 27:72]
  wire  _T_22722 = bht_rd_addr_f == 8'h70; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_112; // @[Reg.scala 27:20]
  wire [1:0] _T_23122 = _T_22722 ? bht_bank_rd_data_out_1_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23377 = _T_23376 | _T_23122; // @[Mux.scala 27:72]
  wire  _T_22724 = bht_rd_addr_f == 8'h71; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_113; // @[Reg.scala 27:20]
  wire [1:0] _T_23123 = _T_22724 ? bht_bank_rd_data_out_1_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23378 = _T_23377 | _T_23123; // @[Mux.scala 27:72]
  wire  _T_22726 = bht_rd_addr_f == 8'h72; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_114; // @[Reg.scala 27:20]
  wire [1:0] _T_23124 = _T_22726 ? bht_bank_rd_data_out_1_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23379 = _T_23378 | _T_23124; // @[Mux.scala 27:72]
  wire  _T_22728 = bht_rd_addr_f == 8'h73; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_115; // @[Reg.scala 27:20]
  wire [1:0] _T_23125 = _T_22728 ? bht_bank_rd_data_out_1_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23380 = _T_23379 | _T_23125; // @[Mux.scala 27:72]
  wire  _T_22730 = bht_rd_addr_f == 8'h74; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_116; // @[Reg.scala 27:20]
  wire [1:0] _T_23126 = _T_22730 ? bht_bank_rd_data_out_1_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23381 = _T_23380 | _T_23126; // @[Mux.scala 27:72]
  wire  _T_22732 = bht_rd_addr_f == 8'h75; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_117; // @[Reg.scala 27:20]
  wire [1:0] _T_23127 = _T_22732 ? bht_bank_rd_data_out_1_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23382 = _T_23381 | _T_23127; // @[Mux.scala 27:72]
  wire  _T_22734 = bht_rd_addr_f == 8'h76; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_118; // @[Reg.scala 27:20]
  wire [1:0] _T_23128 = _T_22734 ? bht_bank_rd_data_out_1_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23383 = _T_23382 | _T_23128; // @[Mux.scala 27:72]
  wire  _T_22736 = bht_rd_addr_f == 8'h77; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_119; // @[Reg.scala 27:20]
  wire [1:0] _T_23129 = _T_22736 ? bht_bank_rd_data_out_1_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23384 = _T_23383 | _T_23129; // @[Mux.scala 27:72]
  wire  _T_22738 = bht_rd_addr_f == 8'h78; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_120; // @[Reg.scala 27:20]
  wire [1:0] _T_23130 = _T_22738 ? bht_bank_rd_data_out_1_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23385 = _T_23384 | _T_23130; // @[Mux.scala 27:72]
  wire  _T_22740 = bht_rd_addr_f == 8'h79; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_121; // @[Reg.scala 27:20]
  wire [1:0] _T_23131 = _T_22740 ? bht_bank_rd_data_out_1_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23386 = _T_23385 | _T_23131; // @[Mux.scala 27:72]
  wire  _T_22742 = bht_rd_addr_f == 8'h7a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_122; // @[Reg.scala 27:20]
  wire [1:0] _T_23132 = _T_22742 ? bht_bank_rd_data_out_1_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23387 = _T_23386 | _T_23132; // @[Mux.scala 27:72]
  wire  _T_22744 = bht_rd_addr_f == 8'h7b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_123; // @[Reg.scala 27:20]
  wire [1:0] _T_23133 = _T_22744 ? bht_bank_rd_data_out_1_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23388 = _T_23387 | _T_23133; // @[Mux.scala 27:72]
  wire  _T_22746 = bht_rd_addr_f == 8'h7c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_124; // @[Reg.scala 27:20]
  wire [1:0] _T_23134 = _T_22746 ? bht_bank_rd_data_out_1_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23389 = _T_23388 | _T_23134; // @[Mux.scala 27:72]
  wire  _T_22748 = bht_rd_addr_f == 8'h7d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_125; // @[Reg.scala 27:20]
  wire [1:0] _T_23135 = _T_22748 ? bht_bank_rd_data_out_1_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23390 = _T_23389 | _T_23135; // @[Mux.scala 27:72]
  wire  _T_22750 = bht_rd_addr_f == 8'h7e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_126; // @[Reg.scala 27:20]
  wire [1:0] _T_23136 = _T_22750 ? bht_bank_rd_data_out_1_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23391 = _T_23390 | _T_23136; // @[Mux.scala 27:72]
  wire  _T_22752 = bht_rd_addr_f == 8'h7f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_127; // @[Reg.scala 27:20]
  wire [1:0] _T_23137 = _T_22752 ? bht_bank_rd_data_out_1_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23392 = _T_23391 | _T_23137; // @[Mux.scala 27:72]
  wire  _T_22754 = bht_rd_addr_f == 8'h80; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_128; // @[Reg.scala 27:20]
  wire [1:0] _T_23138 = _T_22754 ? bht_bank_rd_data_out_1_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23393 = _T_23392 | _T_23138; // @[Mux.scala 27:72]
  wire  _T_22756 = bht_rd_addr_f == 8'h81; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_129; // @[Reg.scala 27:20]
  wire [1:0] _T_23139 = _T_22756 ? bht_bank_rd_data_out_1_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23394 = _T_23393 | _T_23139; // @[Mux.scala 27:72]
  wire  _T_22758 = bht_rd_addr_f == 8'h82; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_130; // @[Reg.scala 27:20]
  wire [1:0] _T_23140 = _T_22758 ? bht_bank_rd_data_out_1_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23395 = _T_23394 | _T_23140; // @[Mux.scala 27:72]
  wire  _T_22760 = bht_rd_addr_f == 8'h83; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_131; // @[Reg.scala 27:20]
  wire [1:0] _T_23141 = _T_22760 ? bht_bank_rd_data_out_1_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23396 = _T_23395 | _T_23141; // @[Mux.scala 27:72]
  wire  _T_22762 = bht_rd_addr_f == 8'h84; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_132; // @[Reg.scala 27:20]
  wire [1:0] _T_23142 = _T_22762 ? bht_bank_rd_data_out_1_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23397 = _T_23396 | _T_23142; // @[Mux.scala 27:72]
  wire  _T_22764 = bht_rd_addr_f == 8'h85; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_133; // @[Reg.scala 27:20]
  wire [1:0] _T_23143 = _T_22764 ? bht_bank_rd_data_out_1_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23398 = _T_23397 | _T_23143; // @[Mux.scala 27:72]
  wire  _T_22766 = bht_rd_addr_f == 8'h86; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_134; // @[Reg.scala 27:20]
  wire [1:0] _T_23144 = _T_22766 ? bht_bank_rd_data_out_1_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23399 = _T_23398 | _T_23144; // @[Mux.scala 27:72]
  wire  _T_22768 = bht_rd_addr_f == 8'h87; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_135; // @[Reg.scala 27:20]
  wire [1:0] _T_23145 = _T_22768 ? bht_bank_rd_data_out_1_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23400 = _T_23399 | _T_23145; // @[Mux.scala 27:72]
  wire  _T_22770 = bht_rd_addr_f == 8'h88; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_136; // @[Reg.scala 27:20]
  wire [1:0] _T_23146 = _T_22770 ? bht_bank_rd_data_out_1_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23401 = _T_23400 | _T_23146; // @[Mux.scala 27:72]
  wire  _T_22772 = bht_rd_addr_f == 8'h89; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_137; // @[Reg.scala 27:20]
  wire [1:0] _T_23147 = _T_22772 ? bht_bank_rd_data_out_1_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23402 = _T_23401 | _T_23147; // @[Mux.scala 27:72]
  wire  _T_22774 = bht_rd_addr_f == 8'h8a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_138; // @[Reg.scala 27:20]
  wire [1:0] _T_23148 = _T_22774 ? bht_bank_rd_data_out_1_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23403 = _T_23402 | _T_23148; // @[Mux.scala 27:72]
  wire  _T_22776 = bht_rd_addr_f == 8'h8b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_139; // @[Reg.scala 27:20]
  wire [1:0] _T_23149 = _T_22776 ? bht_bank_rd_data_out_1_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23404 = _T_23403 | _T_23149; // @[Mux.scala 27:72]
  wire  _T_22778 = bht_rd_addr_f == 8'h8c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_140; // @[Reg.scala 27:20]
  wire [1:0] _T_23150 = _T_22778 ? bht_bank_rd_data_out_1_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23405 = _T_23404 | _T_23150; // @[Mux.scala 27:72]
  wire  _T_22780 = bht_rd_addr_f == 8'h8d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_141; // @[Reg.scala 27:20]
  wire [1:0] _T_23151 = _T_22780 ? bht_bank_rd_data_out_1_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23406 = _T_23405 | _T_23151; // @[Mux.scala 27:72]
  wire  _T_22782 = bht_rd_addr_f == 8'h8e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_142; // @[Reg.scala 27:20]
  wire [1:0] _T_23152 = _T_22782 ? bht_bank_rd_data_out_1_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23407 = _T_23406 | _T_23152; // @[Mux.scala 27:72]
  wire  _T_22784 = bht_rd_addr_f == 8'h8f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_143; // @[Reg.scala 27:20]
  wire [1:0] _T_23153 = _T_22784 ? bht_bank_rd_data_out_1_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23408 = _T_23407 | _T_23153; // @[Mux.scala 27:72]
  wire  _T_22786 = bht_rd_addr_f == 8'h90; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_144; // @[Reg.scala 27:20]
  wire [1:0] _T_23154 = _T_22786 ? bht_bank_rd_data_out_1_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23409 = _T_23408 | _T_23154; // @[Mux.scala 27:72]
  wire  _T_22788 = bht_rd_addr_f == 8'h91; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_145; // @[Reg.scala 27:20]
  wire [1:0] _T_23155 = _T_22788 ? bht_bank_rd_data_out_1_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23410 = _T_23409 | _T_23155; // @[Mux.scala 27:72]
  wire  _T_22790 = bht_rd_addr_f == 8'h92; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_146; // @[Reg.scala 27:20]
  wire [1:0] _T_23156 = _T_22790 ? bht_bank_rd_data_out_1_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23411 = _T_23410 | _T_23156; // @[Mux.scala 27:72]
  wire  _T_22792 = bht_rd_addr_f == 8'h93; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_147; // @[Reg.scala 27:20]
  wire [1:0] _T_23157 = _T_22792 ? bht_bank_rd_data_out_1_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23412 = _T_23411 | _T_23157; // @[Mux.scala 27:72]
  wire  _T_22794 = bht_rd_addr_f == 8'h94; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_148; // @[Reg.scala 27:20]
  wire [1:0] _T_23158 = _T_22794 ? bht_bank_rd_data_out_1_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23413 = _T_23412 | _T_23158; // @[Mux.scala 27:72]
  wire  _T_22796 = bht_rd_addr_f == 8'h95; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_149; // @[Reg.scala 27:20]
  wire [1:0] _T_23159 = _T_22796 ? bht_bank_rd_data_out_1_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23414 = _T_23413 | _T_23159; // @[Mux.scala 27:72]
  wire  _T_22798 = bht_rd_addr_f == 8'h96; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_150; // @[Reg.scala 27:20]
  wire [1:0] _T_23160 = _T_22798 ? bht_bank_rd_data_out_1_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23415 = _T_23414 | _T_23160; // @[Mux.scala 27:72]
  wire  _T_22800 = bht_rd_addr_f == 8'h97; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_151; // @[Reg.scala 27:20]
  wire [1:0] _T_23161 = _T_22800 ? bht_bank_rd_data_out_1_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23416 = _T_23415 | _T_23161; // @[Mux.scala 27:72]
  wire  _T_22802 = bht_rd_addr_f == 8'h98; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_152; // @[Reg.scala 27:20]
  wire [1:0] _T_23162 = _T_22802 ? bht_bank_rd_data_out_1_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23417 = _T_23416 | _T_23162; // @[Mux.scala 27:72]
  wire  _T_22804 = bht_rd_addr_f == 8'h99; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_153; // @[Reg.scala 27:20]
  wire [1:0] _T_23163 = _T_22804 ? bht_bank_rd_data_out_1_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23418 = _T_23417 | _T_23163; // @[Mux.scala 27:72]
  wire  _T_22806 = bht_rd_addr_f == 8'h9a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_154; // @[Reg.scala 27:20]
  wire [1:0] _T_23164 = _T_22806 ? bht_bank_rd_data_out_1_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23419 = _T_23418 | _T_23164; // @[Mux.scala 27:72]
  wire  _T_22808 = bht_rd_addr_f == 8'h9b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_155; // @[Reg.scala 27:20]
  wire [1:0] _T_23165 = _T_22808 ? bht_bank_rd_data_out_1_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23420 = _T_23419 | _T_23165; // @[Mux.scala 27:72]
  wire  _T_22810 = bht_rd_addr_f == 8'h9c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_156; // @[Reg.scala 27:20]
  wire [1:0] _T_23166 = _T_22810 ? bht_bank_rd_data_out_1_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23421 = _T_23420 | _T_23166; // @[Mux.scala 27:72]
  wire  _T_22812 = bht_rd_addr_f == 8'h9d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_157; // @[Reg.scala 27:20]
  wire [1:0] _T_23167 = _T_22812 ? bht_bank_rd_data_out_1_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23422 = _T_23421 | _T_23167; // @[Mux.scala 27:72]
  wire  _T_22814 = bht_rd_addr_f == 8'h9e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_158; // @[Reg.scala 27:20]
  wire [1:0] _T_23168 = _T_22814 ? bht_bank_rd_data_out_1_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23423 = _T_23422 | _T_23168; // @[Mux.scala 27:72]
  wire  _T_22816 = bht_rd_addr_f == 8'h9f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_159; // @[Reg.scala 27:20]
  wire [1:0] _T_23169 = _T_22816 ? bht_bank_rd_data_out_1_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23424 = _T_23423 | _T_23169; // @[Mux.scala 27:72]
  wire  _T_22818 = bht_rd_addr_f == 8'ha0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_160; // @[Reg.scala 27:20]
  wire [1:0] _T_23170 = _T_22818 ? bht_bank_rd_data_out_1_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23425 = _T_23424 | _T_23170; // @[Mux.scala 27:72]
  wire  _T_22820 = bht_rd_addr_f == 8'ha1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_161; // @[Reg.scala 27:20]
  wire [1:0] _T_23171 = _T_22820 ? bht_bank_rd_data_out_1_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23426 = _T_23425 | _T_23171; // @[Mux.scala 27:72]
  wire  _T_22822 = bht_rd_addr_f == 8'ha2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_162; // @[Reg.scala 27:20]
  wire [1:0] _T_23172 = _T_22822 ? bht_bank_rd_data_out_1_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23427 = _T_23426 | _T_23172; // @[Mux.scala 27:72]
  wire  _T_22824 = bht_rd_addr_f == 8'ha3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_163; // @[Reg.scala 27:20]
  wire [1:0] _T_23173 = _T_22824 ? bht_bank_rd_data_out_1_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23428 = _T_23427 | _T_23173; // @[Mux.scala 27:72]
  wire  _T_22826 = bht_rd_addr_f == 8'ha4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_164; // @[Reg.scala 27:20]
  wire [1:0] _T_23174 = _T_22826 ? bht_bank_rd_data_out_1_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23429 = _T_23428 | _T_23174; // @[Mux.scala 27:72]
  wire  _T_22828 = bht_rd_addr_f == 8'ha5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_165; // @[Reg.scala 27:20]
  wire [1:0] _T_23175 = _T_22828 ? bht_bank_rd_data_out_1_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23430 = _T_23429 | _T_23175; // @[Mux.scala 27:72]
  wire  _T_22830 = bht_rd_addr_f == 8'ha6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_166; // @[Reg.scala 27:20]
  wire [1:0] _T_23176 = _T_22830 ? bht_bank_rd_data_out_1_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23431 = _T_23430 | _T_23176; // @[Mux.scala 27:72]
  wire  _T_22832 = bht_rd_addr_f == 8'ha7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_167; // @[Reg.scala 27:20]
  wire [1:0] _T_23177 = _T_22832 ? bht_bank_rd_data_out_1_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23432 = _T_23431 | _T_23177; // @[Mux.scala 27:72]
  wire  _T_22834 = bht_rd_addr_f == 8'ha8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_168; // @[Reg.scala 27:20]
  wire [1:0] _T_23178 = _T_22834 ? bht_bank_rd_data_out_1_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23433 = _T_23432 | _T_23178; // @[Mux.scala 27:72]
  wire  _T_22836 = bht_rd_addr_f == 8'ha9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_169; // @[Reg.scala 27:20]
  wire [1:0] _T_23179 = _T_22836 ? bht_bank_rd_data_out_1_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23434 = _T_23433 | _T_23179; // @[Mux.scala 27:72]
  wire  _T_22838 = bht_rd_addr_f == 8'haa; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_170; // @[Reg.scala 27:20]
  wire [1:0] _T_23180 = _T_22838 ? bht_bank_rd_data_out_1_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23435 = _T_23434 | _T_23180; // @[Mux.scala 27:72]
  wire  _T_22840 = bht_rd_addr_f == 8'hab; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_171; // @[Reg.scala 27:20]
  wire [1:0] _T_23181 = _T_22840 ? bht_bank_rd_data_out_1_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23436 = _T_23435 | _T_23181; // @[Mux.scala 27:72]
  wire  _T_22842 = bht_rd_addr_f == 8'hac; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_172; // @[Reg.scala 27:20]
  wire [1:0] _T_23182 = _T_22842 ? bht_bank_rd_data_out_1_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23437 = _T_23436 | _T_23182; // @[Mux.scala 27:72]
  wire  _T_22844 = bht_rd_addr_f == 8'had; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_173; // @[Reg.scala 27:20]
  wire [1:0] _T_23183 = _T_22844 ? bht_bank_rd_data_out_1_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23438 = _T_23437 | _T_23183; // @[Mux.scala 27:72]
  wire  _T_22846 = bht_rd_addr_f == 8'hae; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_174; // @[Reg.scala 27:20]
  wire [1:0] _T_23184 = _T_22846 ? bht_bank_rd_data_out_1_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23439 = _T_23438 | _T_23184; // @[Mux.scala 27:72]
  wire  _T_22848 = bht_rd_addr_f == 8'haf; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_175; // @[Reg.scala 27:20]
  wire [1:0] _T_23185 = _T_22848 ? bht_bank_rd_data_out_1_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23440 = _T_23439 | _T_23185; // @[Mux.scala 27:72]
  wire  _T_22850 = bht_rd_addr_f == 8'hb0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_176; // @[Reg.scala 27:20]
  wire [1:0] _T_23186 = _T_22850 ? bht_bank_rd_data_out_1_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23441 = _T_23440 | _T_23186; // @[Mux.scala 27:72]
  wire  _T_22852 = bht_rd_addr_f == 8'hb1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_177; // @[Reg.scala 27:20]
  wire [1:0] _T_23187 = _T_22852 ? bht_bank_rd_data_out_1_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23442 = _T_23441 | _T_23187; // @[Mux.scala 27:72]
  wire  _T_22854 = bht_rd_addr_f == 8'hb2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_178; // @[Reg.scala 27:20]
  wire [1:0] _T_23188 = _T_22854 ? bht_bank_rd_data_out_1_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23443 = _T_23442 | _T_23188; // @[Mux.scala 27:72]
  wire  _T_22856 = bht_rd_addr_f == 8'hb3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_179; // @[Reg.scala 27:20]
  wire [1:0] _T_23189 = _T_22856 ? bht_bank_rd_data_out_1_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23444 = _T_23443 | _T_23189; // @[Mux.scala 27:72]
  wire  _T_22858 = bht_rd_addr_f == 8'hb4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_180; // @[Reg.scala 27:20]
  wire [1:0] _T_23190 = _T_22858 ? bht_bank_rd_data_out_1_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23445 = _T_23444 | _T_23190; // @[Mux.scala 27:72]
  wire  _T_22860 = bht_rd_addr_f == 8'hb5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_181; // @[Reg.scala 27:20]
  wire [1:0] _T_23191 = _T_22860 ? bht_bank_rd_data_out_1_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23446 = _T_23445 | _T_23191; // @[Mux.scala 27:72]
  wire  _T_22862 = bht_rd_addr_f == 8'hb6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_182; // @[Reg.scala 27:20]
  wire [1:0] _T_23192 = _T_22862 ? bht_bank_rd_data_out_1_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23447 = _T_23446 | _T_23192; // @[Mux.scala 27:72]
  wire  _T_22864 = bht_rd_addr_f == 8'hb7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_183; // @[Reg.scala 27:20]
  wire [1:0] _T_23193 = _T_22864 ? bht_bank_rd_data_out_1_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23448 = _T_23447 | _T_23193; // @[Mux.scala 27:72]
  wire  _T_22866 = bht_rd_addr_f == 8'hb8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_184; // @[Reg.scala 27:20]
  wire [1:0] _T_23194 = _T_22866 ? bht_bank_rd_data_out_1_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23449 = _T_23448 | _T_23194; // @[Mux.scala 27:72]
  wire  _T_22868 = bht_rd_addr_f == 8'hb9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_185; // @[Reg.scala 27:20]
  wire [1:0] _T_23195 = _T_22868 ? bht_bank_rd_data_out_1_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23450 = _T_23449 | _T_23195; // @[Mux.scala 27:72]
  wire  _T_22870 = bht_rd_addr_f == 8'hba; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_186; // @[Reg.scala 27:20]
  wire [1:0] _T_23196 = _T_22870 ? bht_bank_rd_data_out_1_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23451 = _T_23450 | _T_23196; // @[Mux.scala 27:72]
  wire  _T_22872 = bht_rd_addr_f == 8'hbb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_187; // @[Reg.scala 27:20]
  wire [1:0] _T_23197 = _T_22872 ? bht_bank_rd_data_out_1_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23452 = _T_23451 | _T_23197; // @[Mux.scala 27:72]
  wire  _T_22874 = bht_rd_addr_f == 8'hbc; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_188; // @[Reg.scala 27:20]
  wire [1:0] _T_23198 = _T_22874 ? bht_bank_rd_data_out_1_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23453 = _T_23452 | _T_23198; // @[Mux.scala 27:72]
  wire  _T_22876 = bht_rd_addr_f == 8'hbd; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_189; // @[Reg.scala 27:20]
  wire [1:0] _T_23199 = _T_22876 ? bht_bank_rd_data_out_1_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23454 = _T_23453 | _T_23199; // @[Mux.scala 27:72]
  wire  _T_22878 = bht_rd_addr_f == 8'hbe; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_190; // @[Reg.scala 27:20]
  wire [1:0] _T_23200 = _T_22878 ? bht_bank_rd_data_out_1_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23455 = _T_23454 | _T_23200; // @[Mux.scala 27:72]
  wire  _T_22880 = bht_rd_addr_f == 8'hbf; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_191; // @[Reg.scala 27:20]
  wire [1:0] _T_23201 = _T_22880 ? bht_bank_rd_data_out_1_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23456 = _T_23455 | _T_23201; // @[Mux.scala 27:72]
  wire  _T_22882 = bht_rd_addr_f == 8'hc0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_192; // @[Reg.scala 27:20]
  wire [1:0] _T_23202 = _T_22882 ? bht_bank_rd_data_out_1_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23457 = _T_23456 | _T_23202; // @[Mux.scala 27:72]
  wire  _T_22884 = bht_rd_addr_f == 8'hc1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_193; // @[Reg.scala 27:20]
  wire [1:0] _T_23203 = _T_22884 ? bht_bank_rd_data_out_1_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23458 = _T_23457 | _T_23203; // @[Mux.scala 27:72]
  wire  _T_22886 = bht_rd_addr_f == 8'hc2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_194; // @[Reg.scala 27:20]
  wire [1:0] _T_23204 = _T_22886 ? bht_bank_rd_data_out_1_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23459 = _T_23458 | _T_23204; // @[Mux.scala 27:72]
  wire  _T_22888 = bht_rd_addr_f == 8'hc3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_195; // @[Reg.scala 27:20]
  wire [1:0] _T_23205 = _T_22888 ? bht_bank_rd_data_out_1_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23460 = _T_23459 | _T_23205; // @[Mux.scala 27:72]
  wire  _T_22890 = bht_rd_addr_f == 8'hc4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_196; // @[Reg.scala 27:20]
  wire [1:0] _T_23206 = _T_22890 ? bht_bank_rd_data_out_1_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23461 = _T_23460 | _T_23206; // @[Mux.scala 27:72]
  wire  _T_22892 = bht_rd_addr_f == 8'hc5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_197; // @[Reg.scala 27:20]
  wire [1:0] _T_23207 = _T_22892 ? bht_bank_rd_data_out_1_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23462 = _T_23461 | _T_23207; // @[Mux.scala 27:72]
  wire  _T_22894 = bht_rd_addr_f == 8'hc6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_198; // @[Reg.scala 27:20]
  wire [1:0] _T_23208 = _T_22894 ? bht_bank_rd_data_out_1_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23463 = _T_23462 | _T_23208; // @[Mux.scala 27:72]
  wire  _T_22896 = bht_rd_addr_f == 8'hc7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_199; // @[Reg.scala 27:20]
  wire [1:0] _T_23209 = _T_22896 ? bht_bank_rd_data_out_1_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23464 = _T_23463 | _T_23209; // @[Mux.scala 27:72]
  wire  _T_22898 = bht_rd_addr_f == 8'hc8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_200; // @[Reg.scala 27:20]
  wire [1:0] _T_23210 = _T_22898 ? bht_bank_rd_data_out_1_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23465 = _T_23464 | _T_23210; // @[Mux.scala 27:72]
  wire  _T_22900 = bht_rd_addr_f == 8'hc9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_201; // @[Reg.scala 27:20]
  wire [1:0] _T_23211 = _T_22900 ? bht_bank_rd_data_out_1_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23466 = _T_23465 | _T_23211; // @[Mux.scala 27:72]
  wire  _T_22902 = bht_rd_addr_f == 8'hca; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_202; // @[Reg.scala 27:20]
  wire [1:0] _T_23212 = _T_22902 ? bht_bank_rd_data_out_1_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23467 = _T_23466 | _T_23212; // @[Mux.scala 27:72]
  wire  _T_22904 = bht_rd_addr_f == 8'hcb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_203; // @[Reg.scala 27:20]
  wire [1:0] _T_23213 = _T_22904 ? bht_bank_rd_data_out_1_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23468 = _T_23467 | _T_23213; // @[Mux.scala 27:72]
  wire  _T_22906 = bht_rd_addr_f == 8'hcc; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_204; // @[Reg.scala 27:20]
  wire [1:0] _T_23214 = _T_22906 ? bht_bank_rd_data_out_1_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23469 = _T_23468 | _T_23214; // @[Mux.scala 27:72]
  wire  _T_22908 = bht_rd_addr_f == 8'hcd; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_205; // @[Reg.scala 27:20]
  wire [1:0] _T_23215 = _T_22908 ? bht_bank_rd_data_out_1_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23470 = _T_23469 | _T_23215; // @[Mux.scala 27:72]
  wire  _T_22910 = bht_rd_addr_f == 8'hce; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_206; // @[Reg.scala 27:20]
  wire [1:0] _T_23216 = _T_22910 ? bht_bank_rd_data_out_1_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23471 = _T_23470 | _T_23216; // @[Mux.scala 27:72]
  wire  _T_22912 = bht_rd_addr_f == 8'hcf; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_207; // @[Reg.scala 27:20]
  wire [1:0] _T_23217 = _T_22912 ? bht_bank_rd_data_out_1_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23472 = _T_23471 | _T_23217; // @[Mux.scala 27:72]
  wire  _T_22914 = bht_rd_addr_f == 8'hd0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_208; // @[Reg.scala 27:20]
  wire [1:0] _T_23218 = _T_22914 ? bht_bank_rd_data_out_1_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23473 = _T_23472 | _T_23218; // @[Mux.scala 27:72]
  wire  _T_22916 = bht_rd_addr_f == 8'hd1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_209; // @[Reg.scala 27:20]
  wire [1:0] _T_23219 = _T_22916 ? bht_bank_rd_data_out_1_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23474 = _T_23473 | _T_23219; // @[Mux.scala 27:72]
  wire  _T_22918 = bht_rd_addr_f == 8'hd2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_210; // @[Reg.scala 27:20]
  wire [1:0] _T_23220 = _T_22918 ? bht_bank_rd_data_out_1_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23475 = _T_23474 | _T_23220; // @[Mux.scala 27:72]
  wire  _T_22920 = bht_rd_addr_f == 8'hd3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_211; // @[Reg.scala 27:20]
  wire [1:0] _T_23221 = _T_22920 ? bht_bank_rd_data_out_1_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23476 = _T_23475 | _T_23221; // @[Mux.scala 27:72]
  wire  _T_22922 = bht_rd_addr_f == 8'hd4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_212; // @[Reg.scala 27:20]
  wire [1:0] _T_23222 = _T_22922 ? bht_bank_rd_data_out_1_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23477 = _T_23476 | _T_23222; // @[Mux.scala 27:72]
  wire  _T_22924 = bht_rd_addr_f == 8'hd5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_213; // @[Reg.scala 27:20]
  wire [1:0] _T_23223 = _T_22924 ? bht_bank_rd_data_out_1_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23478 = _T_23477 | _T_23223; // @[Mux.scala 27:72]
  wire  _T_22926 = bht_rd_addr_f == 8'hd6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_214; // @[Reg.scala 27:20]
  wire [1:0] _T_23224 = _T_22926 ? bht_bank_rd_data_out_1_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23479 = _T_23478 | _T_23224; // @[Mux.scala 27:72]
  wire  _T_22928 = bht_rd_addr_f == 8'hd7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_215; // @[Reg.scala 27:20]
  wire [1:0] _T_23225 = _T_22928 ? bht_bank_rd_data_out_1_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23480 = _T_23479 | _T_23225; // @[Mux.scala 27:72]
  wire  _T_22930 = bht_rd_addr_f == 8'hd8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_216; // @[Reg.scala 27:20]
  wire [1:0] _T_23226 = _T_22930 ? bht_bank_rd_data_out_1_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23481 = _T_23480 | _T_23226; // @[Mux.scala 27:72]
  wire  _T_22932 = bht_rd_addr_f == 8'hd9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_217; // @[Reg.scala 27:20]
  wire [1:0] _T_23227 = _T_22932 ? bht_bank_rd_data_out_1_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23482 = _T_23481 | _T_23227; // @[Mux.scala 27:72]
  wire  _T_22934 = bht_rd_addr_f == 8'hda; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_218; // @[Reg.scala 27:20]
  wire [1:0] _T_23228 = _T_22934 ? bht_bank_rd_data_out_1_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23483 = _T_23482 | _T_23228; // @[Mux.scala 27:72]
  wire  _T_22936 = bht_rd_addr_f == 8'hdb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_219; // @[Reg.scala 27:20]
  wire [1:0] _T_23229 = _T_22936 ? bht_bank_rd_data_out_1_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23484 = _T_23483 | _T_23229; // @[Mux.scala 27:72]
  wire  _T_22938 = bht_rd_addr_f == 8'hdc; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_220; // @[Reg.scala 27:20]
  wire [1:0] _T_23230 = _T_22938 ? bht_bank_rd_data_out_1_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23485 = _T_23484 | _T_23230; // @[Mux.scala 27:72]
  wire  _T_22940 = bht_rd_addr_f == 8'hdd; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_221; // @[Reg.scala 27:20]
  wire [1:0] _T_23231 = _T_22940 ? bht_bank_rd_data_out_1_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23486 = _T_23485 | _T_23231; // @[Mux.scala 27:72]
  wire  _T_22942 = bht_rd_addr_f == 8'hde; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_222; // @[Reg.scala 27:20]
  wire [1:0] _T_23232 = _T_22942 ? bht_bank_rd_data_out_1_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23487 = _T_23486 | _T_23232; // @[Mux.scala 27:72]
  wire  _T_22944 = bht_rd_addr_f == 8'hdf; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_223; // @[Reg.scala 27:20]
  wire [1:0] _T_23233 = _T_22944 ? bht_bank_rd_data_out_1_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23488 = _T_23487 | _T_23233; // @[Mux.scala 27:72]
  wire  _T_22946 = bht_rd_addr_f == 8'he0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_224; // @[Reg.scala 27:20]
  wire [1:0] _T_23234 = _T_22946 ? bht_bank_rd_data_out_1_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23489 = _T_23488 | _T_23234; // @[Mux.scala 27:72]
  wire  _T_22948 = bht_rd_addr_f == 8'he1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_225; // @[Reg.scala 27:20]
  wire [1:0] _T_23235 = _T_22948 ? bht_bank_rd_data_out_1_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23490 = _T_23489 | _T_23235; // @[Mux.scala 27:72]
  wire  _T_22950 = bht_rd_addr_f == 8'he2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_226; // @[Reg.scala 27:20]
  wire [1:0] _T_23236 = _T_22950 ? bht_bank_rd_data_out_1_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23491 = _T_23490 | _T_23236; // @[Mux.scala 27:72]
  wire  _T_22952 = bht_rd_addr_f == 8'he3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_227; // @[Reg.scala 27:20]
  wire [1:0] _T_23237 = _T_22952 ? bht_bank_rd_data_out_1_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23492 = _T_23491 | _T_23237; // @[Mux.scala 27:72]
  wire  _T_22954 = bht_rd_addr_f == 8'he4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_228; // @[Reg.scala 27:20]
  wire [1:0] _T_23238 = _T_22954 ? bht_bank_rd_data_out_1_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23493 = _T_23492 | _T_23238; // @[Mux.scala 27:72]
  wire  _T_22956 = bht_rd_addr_f == 8'he5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_229; // @[Reg.scala 27:20]
  wire [1:0] _T_23239 = _T_22956 ? bht_bank_rd_data_out_1_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23494 = _T_23493 | _T_23239; // @[Mux.scala 27:72]
  wire  _T_22958 = bht_rd_addr_f == 8'he6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_230; // @[Reg.scala 27:20]
  wire [1:0] _T_23240 = _T_22958 ? bht_bank_rd_data_out_1_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23495 = _T_23494 | _T_23240; // @[Mux.scala 27:72]
  wire  _T_22960 = bht_rd_addr_f == 8'he7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_231; // @[Reg.scala 27:20]
  wire [1:0] _T_23241 = _T_22960 ? bht_bank_rd_data_out_1_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23496 = _T_23495 | _T_23241; // @[Mux.scala 27:72]
  wire  _T_22962 = bht_rd_addr_f == 8'he8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_232; // @[Reg.scala 27:20]
  wire [1:0] _T_23242 = _T_22962 ? bht_bank_rd_data_out_1_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23497 = _T_23496 | _T_23242; // @[Mux.scala 27:72]
  wire  _T_22964 = bht_rd_addr_f == 8'he9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_233; // @[Reg.scala 27:20]
  wire [1:0] _T_23243 = _T_22964 ? bht_bank_rd_data_out_1_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23498 = _T_23497 | _T_23243; // @[Mux.scala 27:72]
  wire  _T_22966 = bht_rd_addr_f == 8'hea; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_234; // @[Reg.scala 27:20]
  wire [1:0] _T_23244 = _T_22966 ? bht_bank_rd_data_out_1_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23499 = _T_23498 | _T_23244; // @[Mux.scala 27:72]
  wire  _T_22968 = bht_rd_addr_f == 8'heb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_235; // @[Reg.scala 27:20]
  wire [1:0] _T_23245 = _T_22968 ? bht_bank_rd_data_out_1_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23500 = _T_23499 | _T_23245; // @[Mux.scala 27:72]
  wire  _T_22970 = bht_rd_addr_f == 8'hec; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_236; // @[Reg.scala 27:20]
  wire [1:0] _T_23246 = _T_22970 ? bht_bank_rd_data_out_1_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23501 = _T_23500 | _T_23246; // @[Mux.scala 27:72]
  wire  _T_22972 = bht_rd_addr_f == 8'hed; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_237; // @[Reg.scala 27:20]
  wire [1:0] _T_23247 = _T_22972 ? bht_bank_rd_data_out_1_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23502 = _T_23501 | _T_23247; // @[Mux.scala 27:72]
  wire  _T_22974 = bht_rd_addr_f == 8'hee; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_238; // @[Reg.scala 27:20]
  wire [1:0] _T_23248 = _T_22974 ? bht_bank_rd_data_out_1_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23503 = _T_23502 | _T_23248; // @[Mux.scala 27:72]
  wire  _T_22976 = bht_rd_addr_f == 8'hef; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_239; // @[Reg.scala 27:20]
  wire [1:0] _T_23249 = _T_22976 ? bht_bank_rd_data_out_1_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23504 = _T_23503 | _T_23249; // @[Mux.scala 27:72]
  wire  _T_22978 = bht_rd_addr_f == 8'hf0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_240; // @[Reg.scala 27:20]
  wire [1:0] _T_23250 = _T_22978 ? bht_bank_rd_data_out_1_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23505 = _T_23504 | _T_23250; // @[Mux.scala 27:72]
  wire  _T_22980 = bht_rd_addr_f == 8'hf1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_241; // @[Reg.scala 27:20]
  wire [1:0] _T_23251 = _T_22980 ? bht_bank_rd_data_out_1_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23506 = _T_23505 | _T_23251; // @[Mux.scala 27:72]
  wire  _T_22982 = bht_rd_addr_f == 8'hf2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_242; // @[Reg.scala 27:20]
  wire [1:0] _T_23252 = _T_22982 ? bht_bank_rd_data_out_1_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23507 = _T_23506 | _T_23252; // @[Mux.scala 27:72]
  wire  _T_22984 = bht_rd_addr_f == 8'hf3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_243; // @[Reg.scala 27:20]
  wire [1:0] _T_23253 = _T_22984 ? bht_bank_rd_data_out_1_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23508 = _T_23507 | _T_23253; // @[Mux.scala 27:72]
  wire  _T_22986 = bht_rd_addr_f == 8'hf4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_244; // @[Reg.scala 27:20]
  wire [1:0] _T_23254 = _T_22986 ? bht_bank_rd_data_out_1_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23509 = _T_23508 | _T_23254; // @[Mux.scala 27:72]
  wire  _T_22988 = bht_rd_addr_f == 8'hf5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_245; // @[Reg.scala 27:20]
  wire [1:0] _T_23255 = _T_22988 ? bht_bank_rd_data_out_1_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23510 = _T_23509 | _T_23255; // @[Mux.scala 27:72]
  wire  _T_22990 = bht_rd_addr_f == 8'hf6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_246; // @[Reg.scala 27:20]
  wire [1:0] _T_23256 = _T_22990 ? bht_bank_rd_data_out_1_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23511 = _T_23510 | _T_23256; // @[Mux.scala 27:72]
  wire  _T_22992 = bht_rd_addr_f == 8'hf7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_247; // @[Reg.scala 27:20]
  wire [1:0] _T_23257 = _T_22992 ? bht_bank_rd_data_out_1_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23512 = _T_23511 | _T_23257; // @[Mux.scala 27:72]
  wire  _T_22994 = bht_rd_addr_f == 8'hf8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_248; // @[Reg.scala 27:20]
  wire [1:0] _T_23258 = _T_22994 ? bht_bank_rd_data_out_1_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23513 = _T_23512 | _T_23258; // @[Mux.scala 27:72]
  wire  _T_22996 = bht_rd_addr_f == 8'hf9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_249; // @[Reg.scala 27:20]
  wire [1:0] _T_23259 = _T_22996 ? bht_bank_rd_data_out_1_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23514 = _T_23513 | _T_23259; // @[Mux.scala 27:72]
  wire  _T_22998 = bht_rd_addr_f == 8'hfa; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_250; // @[Reg.scala 27:20]
  wire [1:0] _T_23260 = _T_22998 ? bht_bank_rd_data_out_1_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23515 = _T_23514 | _T_23260; // @[Mux.scala 27:72]
  wire  _T_23000 = bht_rd_addr_f == 8'hfb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_251; // @[Reg.scala 27:20]
  wire [1:0] _T_23261 = _T_23000 ? bht_bank_rd_data_out_1_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23516 = _T_23515 | _T_23261; // @[Mux.scala 27:72]
  wire  _T_23002 = bht_rd_addr_f == 8'hfc; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_252; // @[Reg.scala 27:20]
  wire [1:0] _T_23262 = _T_23002 ? bht_bank_rd_data_out_1_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23517 = _T_23516 | _T_23262; // @[Mux.scala 27:72]
  wire  _T_23004 = bht_rd_addr_f == 8'hfd; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_253; // @[Reg.scala 27:20]
  wire [1:0] _T_23263 = _T_23004 ? bht_bank_rd_data_out_1_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23518 = _T_23517 | _T_23263; // @[Mux.scala 27:72]
  wire  _T_23006 = bht_rd_addr_f == 8'hfe; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_254; // @[Reg.scala 27:20]
  wire [1:0] _T_23264 = _T_23006 ? bht_bank_rd_data_out_1_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23519 = _T_23518 | _T_23264; // @[Mux.scala 27:72]
  wire  _T_23008 = bht_rd_addr_f == 8'hff; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_255; // @[Reg.scala 27:20]
  wire [1:0] _T_23265 = _T_23008 ? bht_bank_rd_data_out_1_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank1_rd_data_f = _T_23519 | _T_23265; // @[Mux.scala 27:72]
  wire [1:0] _T_279 = _T_162 ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [9:0] _T_611 = {btb_rd_addr_p1_f,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_rd_addr_hashed_p1_f = _T_611[9:2] ^ fghr; // @[lib.scala 56:35]
  wire  _T_23522 = bht_rd_addr_hashed_p1_f == 8'h0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_0; // @[Reg.scala 27:20]
  wire [1:0] _T_24034 = _T_23522 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_23524 = bht_rd_addr_hashed_p1_f == 8'h1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_1; // @[Reg.scala 27:20]
  wire [1:0] _T_24035 = _T_23524 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24290 = _T_24034 | _T_24035; // @[Mux.scala 27:72]
  wire  _T_23526 = bht_rd_addr_hashed_p1_f == 8'h2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_2; // @[Reg.scala 27:20]
  wire [1:0] _T_24036 = _T_23526 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24291 = _T_24290 | _T_24036; // @[Mux.scala 27:72]
  wire  _T_23528 = bht_rd_addr_hashed_p1_f == 8'h3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_3; // @[Reg.scala 27:20]
  wire [1:0] _T_24037 = _T_23528 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24292 = _T_24291 | _T_24037; // @[Mux.scala 27:72]
  wire  _T_23530 = bht_rd_addr_hashed_p1_f == 8'h4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_4; // @[Reg.scala 27:20]
  wire [1:0] _T_24038 = _T_23530 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24293 = _T_24292 | _T_24038; // @[Mux.scala 27:72]
  wire  _T_23532 = bht_rd_addr_hashed_p1_f == 8'h5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_5; // @[Reg.scala 27:20]
  wire [1:0] _T_24039 = _T_23532 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24294 = _T_24293 | _T_24039; // @[Mux.scala 27:72]
  wire  _T_23534 = bht_rd_addr_hashed_p1_f == 8'h6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_6; // @[Reg.scala 27:20]
  wire [1:0] _T_24040 = _T_23534 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24295 = _T_24294 | _T_24040; // @[Mux.scala 27:72]
  wire  _T_23536 = bht_rd_addr_hashed_p1_f == 8'h7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_7; // @[Reg.scala 27:20]
  wire [1:0] _T_24041 = _T_23536 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24296 = _T_24295 | _T_24041; // @[Mux.scala 27:72]
  wire  _T_23538 = bht_rd_addr_hashed_p1_f == 8'h8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_8; // @[Reg.scala 27:20]
  wire [1:0] _T_24042 = _T_23538 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24297 = _T_24296 | _T_24042; // @[Mux.scala 27:72]
  wire  _T_23540 = bht_rd_addr_hashed_p1_f == 8'h9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_9; // @[Reg.scala 27:20]
  wire [1:0] _T_24043 = _T_23540 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24298 = _T_24297 | _T_24043; // @[Mux.scala 27:72]
  wire  _T_23542 = bht_rd_addr_hashed_p1_f == 8'ha; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_10; // @[Reg.scala 27:20]
  wire [1:0] _T_24044 = _T_23542 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24299 = _T_24298 | _T_24044; // @[Mux.scala 27:72]
  wire  _T_23544 = bht_rd_addr_hashed_p1_f == 8'hb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_11; // @[Reg.scala 27:20]
  wire [1:0] _T_24045 = _T_23544 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24300 = _T_24299 | _T_24045; // @[Mux.scala 27:72]
  wire  _T_23546 = bht_rd_addr_hashed_p1_f == 8'hc; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_12; // @[Reg.scala 27:20]
  wire [1:0] _T_24046 = _T_23546 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24301 = _T_24300 | _T_24046; // @[Mux.scala 27:72]
  wire  _T_23548 = bht_rd_addr_hashed_p1_f == 8'hd; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_13; // @[Reg.scala 27:20]
  wire [1:0] _T_24047 = _T_23548 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24302 = _T_24301 | _T_24047; // @[Mux.scala 27:72]
  wire  _T_23550 = bht_rd_addr_hashed_p1_f == 8'he; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_14; // @[Reg.scala 27:20]
  wire [1:0] _T_24048 = _T_23550 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24303 = _T_24302 | _T_24048; // @[Mux.scala 27:72]
  wire  _T_23552 = bht_rd_addr_hashed_p1_f == 8'hf; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_15; // @[Reg.scala 27:20]
  wire [1:0] _T_24049 = _T_23552 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24304 = _T_24303 | _T_24049; // @[Mux.scala 27:72]
  wire  _T_23554 = bht_rd_addr_hashed_p1_f == 8'h10; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_16; // @[Reg.scala 27:20]
  wire [1:0] _T_24050 = _T_23554 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24305 = _T_24304 | _T_24050; // @[Mux.scala 27:72]
  wire  _T_23556 = bht_rd_addr_hashed_p1_f == 8'h11; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_17; // @[Reg.scala 27:20]
  wire [1:0] _T_24051 = _T_23556 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24306 = _T_24305 | _T_24051; // @[Mux.scala 27:72]
  wire  _T_23558 = bht_rd_addr_hashed_p1_f == 8'h12; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_18; // @[Reg.scala 27:20]
  wire [1:0] _T_24052 = _T_23558 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24307 = _T_24306 | _T_24052; // @[Mux.scala 27:72]
  wire  _T_23560 = bht_rd_addr_hashed_p1_f == 8'h13; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_19; // @[Reg.scala 27:20]
  wire [1:0] _T_24053 = _T_23560 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24308 = _T_24307 | _T_24053; // @[Mux.scala 27:72]
  wire  _T_23562 = bht_rd_addr_hashed_p1_f == 8'h14; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_20; // @[Reg.scala 27:20]
  wire [1:0] _T_24054 = _T_23562 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24309 = _T_24308 | _T_24054; // @[Mux.scala 27:72]
  wire  _T_23564 = bht_rd_addr_hashed_p1_f == 8'h15; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_21; // @[Reg.scala 27:20]
  wire [1:0] _T_24055 = _T_23564 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24310 = _T_24309 | _T_24055; // @[Mux.scala 27:72]
  wire  _T_23566 = bht_rd_addr_hashed_p1_f == 8'h16; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_22; // @[Reg.scala 27:20]
  wire [1:0] _T_24056 = _T_23566 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24311 = _T_24310 | _T_24056; // @[Mux.scala 27:72]
  wire  _T_23568 = bht_rd_addr_hashed_p1_f == 8'h17; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_23; // @[Reg.scala 27:20]
  wire [1:0] _T_24057 = _T_23568 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24312 = _T_24311 | _T_24057; // @[Mux.scala 27:72]
  wire  _T_23570 = bht_rd_addr_hashed_p1_f == 8'h18; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_24; // @[Reg.scala 27:20]
  wire [1:0] _T_24058 = _T_23570 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24313 = _T_24312 | _T_24058; // @[Mux.scala 27:72]
  wire  _T_23572 = bht_rd_addr_hashed_p1_f == 8'h19; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_25; // @[Reg.scala 27:20]
  wire [1:0] _T_24059 = _T_23572 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24314 = _T_24313 | _T_24059; // @[Mux.scala 27:72]
  wire  _T_23574 = bht_rd_addr_hashed_p1_f == 8'h1a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_26; // @[Reg.scala 27:20]
  wire [1:0] _T_24060 = _T_23574 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24315 = _T_24314 | _T_24060; // @[Mux.scala 27:72]
  wire  _T_23576 = bht_rd_addr_hashed_p1_f == 8'h1b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_27; // @[Reg.scala 27:20]
  wire [1:0] _T_24061 = _T_23576 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24316 = _T_24315 | _T_24061; // @[Mux.scala 27:72]
  wire  _T_23578 = bht_rd_addr_hashed_p1_f == 8'h1c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_28; // @[Reg.scala 27:20]
  wire [1:0] _T_24062 = _T_23578 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24317 = _T_24316 | _T_24062; // @[Mux.scala 27:72]
  wire  _T_23580 = bht_rd_addr_hashed_p1_f == 8'h1d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_29; // @[Reg.scala 27:20]
  wire [1:0] _T_24063 = _T_23580 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24318 = _T_24317 | _T_24063; // @[Mux.scala 27:72]
  wire  _T_23582 = bht_rd_addr_hashed_p1_f == 8'h1e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_30; // @[Reg.scala 27:20]
  wire [1:0] _T_24064 = _T_23582 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24319 = _T_24318 | _T_24064; // @[Mux.scala 27:72]
  wire  _T_23584 = bht_rd_addr_hashed_p1_f == 8'h1f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_31; // @[Reg.scala 27:20]
  wire [1:0] _T_24065 = _T_23584 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24320 = _T_24319 | _T_24065; // @[Mux.scala 27:72]
  wire  _T_23586 = bht_rd_addr_hashed_p1_f == 8'h20; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_32; // @[Reg.scala 27:20]
  wire [1:0] _T_24066 = _T_23586 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24321 = _T_24320 | _T_24066; // @[Mux.scala 27:72]
  wire  _T_23588 = bht_rd_addr_hashed_p1_f == 8'h21; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_33; // @[Reg.scala 27:20]
  wire [1:0] _T_24067 = _T_23588 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24322 = _T_24321 | _T_24067; // @[Mux.scala 27:72]
  wire  _T_23590 = bht_rd_addr_hashed_p1_f == 8'h22; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_34; // @[Reg.scala 27:20]
  wire [1:0] _T_24068 = _T_23590 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24323 = _T_24322 | _T_24068; // @[Mux.scala 27:72]
  wire  _T_23592 = bht_rd_addr_hashed_p1_f == 8'h23; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_35; // @[Reg.scala 27:20]
  wire [1:0] _T_24069 = _T_23592 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24324 = _T_24323 | _T_24069; // @[Mux.scala 27:72]
  wire  _T_23594 = bht_rd_addr_hashed_p1_f == 8'h24; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_36; // @[Reg.scala 27:20]
  wire [1:0] _T_24070 = _T_23594 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24325 = _T_24324 | _T_24070; // @[Mux.scala 27:72]
  wire  _T_23596 = bht_rd_addr_hashed_p1_f == 8'h25; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_37; // @[Reg.scala 27:20]
  wire [1:0] _T_24071 = _T_23596 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24326 = _T_24325 | _T_24071; // @[Mux.scala 27:72]
  wire  _T_23598 = bht_rd_addr_hashed_p1_f == 8'h26; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_38; // @[Reg.scala 27:20]
  wire [1:0] _T_24072 = _T_23598 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24327 = _T_24326 | _T_24072; // @[Mux.scala 27:72]
  wire  _T_23600 = bht_rd_addr_hashed_p1_f == 8'h27; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_39; // @[Reg.scala 27:20]
  wire [1:0] _T_24073 = _T_23600 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24328 = _T_24327 | _T_24073; // @[Mux.scala 27:72]
  wire  _T_23602 = bht_rd_addr_hashed_p1_f == 8'h28; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_40; // @[Reg.scala 27:20]
  wire [1:0] _T_24074 = _T_23602 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24329 = _T_24328 | _T_24074; // @[Mux.scala 27:72]
  wire  _T_23604 = bht_rd_addr_hashed_p1_f == 8'h29; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_41; // @[Reg.scala 27:20]
  wire [1:0] _T_24075 = _T_23604 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24330 = _T_24329 | _T_24075; // @[Mux.scala 27:72]
  wire  _T_23606 = bht_rd_addr_hashed_p1_f == 8'h2a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_42; // @[Reg.scala 27:20]
  wire [1:0] _T_24076 = _T_23606 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24331 = _T_24330 | _T_24076; // @[Mux.scala 27:72]
  wire  _T_23608 = bht_rd_addr_hashed_p1_f == 8'h2b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_43; // @[Reg.scala 27:20]
  wire [1:0] _T_24077 = _T_23608 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24332 = _T_24331 | _T_24077; // @[Mux.scala 27:72]
  wire  _T_23610 = bht_rd_addr_hashed_p1_f == 8'h2c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_44; // @[Reg.scala 27:20]
  wire [1:0] _T_24078 = _T_23610 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24333 = _T_24332 | _T_24078; // @[Mux.scala 27:72]
  wire  _T_23612 = bht_rd_addr_hashed_p1_f == 8'h2d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_45; // @[Reg.scala 27:20]
  wire [1:0] _T_24079 = _T_23612 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24334 = _T_24333 | _T_24079; // @[Mux.scala 27:72]
  wire  _T_23614 = bht_rd_addr_hashed_p1_f == 8'h2e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_46; // @[Reg.scala 27:20]
  wire [1:0] _T_24080 = _T_23614 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24335 = _T_24334 | _T_24080; // @[Mux.scala 27:72]
  wire  _T_23616 = bht_rd_addr_hashed_p1_f == 8'h2f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_47; // @[Reg.scala 27:20]
  wire [1:0] _T_24081 = _T_23616 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24336 = _T_24335 | _T_24081; // @[Mux.scala 27:72]
  wire  _T_23618 = bht_rd_addr_hashed_p1_f == 8'h30; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_48; // @[Reg.scala 27:20]
  wire [1:0] _T_24082 = _T_23618 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24337 = _T_24336 | _T_24082; // @[Mux.scala 27:72]
  wire  _T_23620 = bht_rd_addr_hashed_p1_f == 8'h31; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_49; // @[Reg.scala 27:20]
  wire [1:0] _T_24083 = _T_23620 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24338 = _T_24337 | _T_24083; // @[Mux.scala 27:72]
  wire  _T_23622 = bht_rd_addr_hashed_p1_f == 8'h32; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_50; // @[Reg.scala 27:20]
  wire [1:0] _T_24084 = _T_23622 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24339 = _T_24338 | _T_24084; // @[Mux.scala 27:72]
  wire  _T_23624 = bht_rd_addr_hashed_p1_f == 8'h33; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_51; // @[Reg.scala 27:20]
  wire [1:0] _T_24085 = _T_23624 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24340 = _T_24339 | _T_24085; // @[Mux.scala 27:72]
  wire  _T_23626 = bht_rd_addr_hashed_p1_f == 8'h34; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_52; // @[Reg.scala 27:20]
  wire [1:0] _T_24086 = _T_23626 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24341 = _T_24340 | _T_24086; // @[Mux.scala 27:72]
  wire  _T_23628 = bht_rd_addr_hashed_p1_f == 8'h35; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_53; // @[Reg.scala 27:20]
  wire [1:0] _T_24087 = _T_23628 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24342 = _T_24341 | _T_24087; // @[Mux.scala 27:72]
  wire  _T_23630 = bht_rd_addr_hashed_p1_f == 8'h36; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_54; // @[Reg.scala 27:20]
  wire [1:0] _T_24088 = _T_23630 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24343 = _T_24342 | _T_24088; // @[Mux.scala 27:72]
  wire  _T_23632 = bht_rd_addr_hashed_p1_f == 8'h37; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_55; // @[Reg.scala 27:20]
  wire [1:0] _T_24089 = _T_23632 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24344 = _T_24343 | _T_24089; // @[Mux.scala 27:72]
  wire  _T_23634 = bht_rd_addr_hashed_p1_f == 8'h38; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_56; // @[Reg.scala 27:20]
  wire [1:0] _T_24090 = _T_23634 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24345 = _T_24344 | _T_24090; // @[Mux.scala 27:72]
  wire  _T_23636 = bht_rd_addr_hashed_p1_f == 8'h39; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_57; // @[Reg.scala 27:20]
  wire [1:0] _T_24091 = _T_23636 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24346 = _T_24345 | _T_24091; // @[Mux.scala 27:72]
  wire  _T_23638 = bht_rd_addr_hashed_p1_f == 8'h3a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_58; // @[Reg.scala 27:20]
  wire [1:0] _T_24092 = _T_23638 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24347 = _T_24346 | _T_24092; // @[Mux.scala 27:72]
  wire  _T_23640 = bht_rd_addr_hashed_p1_f == 8'h3b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_59; // @[Reg.scala 27:20]
  wire [1:0] _T_24093 = _T_23640 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24348 = _T_24347 | _T_24093; // @[Mux.scala 27:72]
  wire  _T_23642 = bht_rd_addr_hashed_p1_f == 8'h3c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_60; // @[Reg.scala 27:20]
  wire [1:0] _T_24094 = _T_23642 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24349 = _T_24348 | _T_24094; // @[Mux.scala 27:72]
  wire  _T_23644 = bht_rd_addr_hashed_p1_f == 8'h3d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_61; // @[Reg.scala 27:20]
  wire [1:0] _T_24095 = _T_23644 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24350 = _T_24349 | _T_24095; // @[Mux.scala 27:72]
  wire  _T_23646 = bht_rd_addr_hashed_p1_f == 8'h3e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_62; // @[Reg.scala 27:20]
  wire [1:0] _T_24096 = _T_23646 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24351 = _T_24350 | _T_24096; // @[Mux.scala 27:72]
  wire  _T_23648 = bht_rd_addr_hashed_p1_f == 8'h3f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_63; // @[Reg.scala 27:20]
  wire [1:0] _T_24097 = _T_23648 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24352 = _T_24351 | _T_24097; // @[Mux.scala 27:72]
  wire  _T_23650 = bht_rd_addr_hashed_p1_f == 8'h40; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_64; // @[Reg.scala 27:20]
  wire [1:0] _T_24098 = _T_23650 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24353 = _T_24352 | _T_24098; // @[Mux.scala 27:72]
  wire  _T_23652 = bht_rd_addr_hashed_p1_f == 8'h41; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_65; // @[Reg.scala 27:20]
  wire [1:0] _T_24099 = _T_23652 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24354 = _T_24353 | _T_24099; // @[Mux.scala 27:72]
  wire  _T_23654 = bht_rd_addr_hashed_p1_f == 8'h42; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_66; // @[Reg.scala 27:20]
  wire [1:0] _T_24100 = _T_23654 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24355 = _T_24354 | _T_24100; // @[Mux.scala 27:72]
  wire  _T_23656 = bht_rd_addr_hashed_p1_f == 8'h43; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_67; // @[Reg.scala 27:20]
  wire [1:0] _T_24101 = _T_23656 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24356 = _T_24355 | _T_24101; // @[Mux.scala 27:72]
  wire  _T_23658 = bht_rd_addr_hashed_p1_f == 8'h44; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_68; // @[Reg.scala 27:20]
  wire [1:0] _T_24102 = _T_23658 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24357 = _T_24356 | _T_24102; // @[Mux.scala 27:72]
  wire  _T_23660 = bht_rd_addr_hashed_p1_f == 8'h45; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_69; // @[Reg.scala 27:20]
  wire [1:0] _T_24103 = _T_23660 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24358 = _T_24357 | _T_24103; // @[Mux.scala 27:72]
  wire  _T_23662 = bht_rd_addr_hashed_p1_f == 8'h46; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_70; // @[Reg.scala 27:20]
  wire [1:0] _T_24104 = _T_23662 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24359 = _T_24358 | _T_24104; // @[Mux.scala 27:72]
  wire  _T_23664 = bht_rd_addr_hashed_p1_f == 8'h47; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_71; // @[Reg.scala 27:20]
  wire [1:0] _T_24105 = _T_23664 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24360 = _T_24359 | _T_24105; // @[Mux.scala 27:72]
  wire  _T_23666 = bht_rd_addr_hashed_p1_f == 8'h48; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_72; // @[Reg.scala 27:20]
  wire [1:0] _T_24106 = _T_23666 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24361 = _T_24360 | _T_24106; // @[Mux.scala 27:72]
  wire  _T_23668 = bht_rd_addr_hashed_p1_f == 8'h49; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_73; // @[Reg.scala 27:20]
  wire [1:0] _T_24107 = _T_23668 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24362 = _T_24361 | _T_24107; // @[Mux.scala 27:72]
  wire  _T_23670 = bht_rd_addr_hashed_p1_f == 8'h4a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_74; // @[Reg.scala 27:20]
  wire [1:0] _T_24108 = _T_23670 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24363 = _T_24362 | _T_24108; // @[Mux.scala 27:72]
  wire  _T_23672 = bht_rd_addr_hashed_p1_f == 8'h4b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_75; // @[Reg.scala 27:20]
  wire [1:0] _T_24109 = _T_23672 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24364 = _T_24363 | _T_24109; // @[Mux.scala 27:72]
  wire  _T_23674 = bht_rd_addr_hashed_p1_f == 8'h4c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_76; // @[Reg.scala 27:20]
  wire [1:0] _T_24110 = _T_23674 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24365 = _T_24364 | _T_24110; // @[Mux.scala 27:72]
  wire  _T_23676 = bht_rd_addr_hashed_p1_f == 8'h4d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_77; // @[Reg.scala 27:20]
  wire [1:0] _T_24111 = _T_23676 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24366 = _T_24365 | _T_24111; // @[Mux.scala 27:72]
  wire  _T_23678 = bht_rd_addr_hashed_p1_f == 8'h4e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_78; // @[Reg.scala 27:20]
  wire [1:0] _T_24112 = _T_23678 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24367 = _T_24366 | _T_24112; // @[Mux.scala 27:72]
  wire  _T_23680 = bht_rd_addr_hashed_p1_f == 8'h4f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_79; // @[Reg.scala 27:20]
  wire [1:0] _T_24113 = _T_23680 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24368 = _T_24367 | _T_24113; // @[Mux.scala 27:72]
  wire  _T_23682 = bht_rd_addr_hashed_p1_f == 8'h50; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_80; // @[Reg.scala 27:20]
  wire [1:0] _T_24114 = _T_23682 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24369 = _T_24368 | _T_24114; // @[Mux.scala 27:72]
  wire  _T_23684 = bht_rd_addr_hashed_p1_f == 8'h51; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_81; // @[Reg.scala 27:20]
  wire [1:0] _T_24115 = _T_23684 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24370 = _T_24369 | _T_24115; // @[Mux.scala 27:72]
  wire  _T_23686 = bht_rd_addr_hashed_p1_f == 8'h52; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_82; // @[Reg.scala 27:20]
  wire [1:0] _T_24116 = _T_23686 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24371 = _T_24370 | _T_24116; // @[Mux.scala 27:72]
  wire  _T_23688 = bht_rd_addr_hashed_p1_f == 8'h53; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_83; // @[Reg.scala 27:20]
  wire [1:0] _T_24117 = _T_23688 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24372 = _T_24371 | _T_24117; // @[Mux.scala 27:72]
  wire  _T_23690 = bht_rd_addr_hashed_p1_f == 8'h54; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_84; // @[Reg.scala 27:20]
  wire [1:0] _T_24118 = _T_23690 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24373 = _T_24372 | _T_24118; // @[Mux.scala 27:72]
  wire  _T_23692 = bht_rd_addr_hashed_p1_f == 8'h55; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_85; // @[Reg.scala 27:20]
  wire [1:0] _T_24119 = _T_23692 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24374 = _T_24373 | _T_24119; // @[Mux.scala 27:72]
  wire  _T_23694 = bht_rd_addr_hashed_p1_f == 8'h56; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_86; // @[Reg.scala 27:20]
  wire [1:0] _T_24120 = _T_23694 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24375 = _T_24374 | _T_24120; // @[Mux.scala 27:72]
  wire  _T_23696 = bht_rd_addr_hashed_p1_f == 8'h57; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_87; // @[Reg.scala 27:20]
  wire [1:0] _T_24121 = _T_23696 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24376 = _T_24375 | _T_24121; // @[Mux.scala 27:72]
  wire  _T_23698 = bht_rd_addr_hashed_p1_f == 8'h58; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_88; // @[Reg.scala 27:20]
  wire [1:0] _T_24122 = _T_23698 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24377 = _T_24376 | _T_24122; // @[Mux.scala 27:72]
  wire  _T_23700 = bht_rd_addr_hashed_p1_f == 8'h59; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_89; // @[Reg.scala 27:20]
  wire [1:0] _T_24123 = _T_23700 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24378 = _T_24377 | _T_24123; // @[Mux.scala 27:72]
  wire  _T_23702 = bht_rd_addr_hashed_p1_f == 8'h5a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_90; // @[Reg.scala 27:20]
  wire [1:0] _T_24124 = _T_23702 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24379 = _T_24378 | _T_24124; // @[Mux.scala 27:72]
  wire  _T_23704 = bht_rd_addr_hashed_p1_f == 8'h5b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_91; // @[Reg.scala 27:20]
  wire [1:0] _T_24125 = _T_23704 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24380 = _T_24379 | _T_24125; // @[Mux.scala 27:72]
  wire  _T_23706 = bht_rd_addr_hashed_p1_f == 8'h5c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_92; // @[Reg.scala 27:20]
  wire [1:0] _T_24126 = _T_23706 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24381 = _T_24380 | _T_24126; // @[Mux.scala 27:72]
  wire  _T_23708 = bht_rd_addr_hashed_p1_f == 8'h5d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_93; // @[Reg.scala 27:20]
  wire [1:0] _T_24127 = _T_23708 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24382 = _T_24381 | _T_24127; // @[Mux.scala 27:72]
  wire  _T_23710 = bht_rd_addr_hashed_p1_f == 8'h5e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_94; // @[Reg.scala 27:20]
  wire [1:0] _T_24128 = _T_23710 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24383 = _T_24382 | _T_24128; // @[Mux.scala 27:72]
  wire  _T_23712 = bht_rd_addr_hashed_p1_f == 8'h5f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_95; // @[Reg.scala 27:20]
  wire [1:0] _T_24129 = _T_23712 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24384 = _T_24383 | _T_24129; // @[Mux.scala 27:72]
  wire  _T_23714 = bht_rd_addr_hashed_p1_f == 8'h60; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_96; // @[Reg.scala 27:20]
  wire [1:0] _T_24130 = _T_23714 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24385 = _T_24384 | _T_24130; // @[Mux.scala 27:72]
  wire  _T_23716 = bht_rd_addr_hashed_p1_f == 8'h61; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_97; // @[Reg.scala 27:20]
  wire [1:0] _T_24131 = _T_23716 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24386 = _T_24385 | _T_24131; // @[Mux.scala 27:72]
  wire  _T_23718 = bht_rd_addr_hashed_p1_f == 8'h62; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_98; // @[Reg.scala 27:20]
  wire [1:0] _T_24132 = _T_23718 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24387 = _T_24386 | _T_24132; // @[Mux.scala 27:72]
  wire  _T_23720 = bht_rd_addr_hashed_p1_f == 8'h63; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_99; // @[Reg.scala 27:20]
  wire [1:0] _T_24133 = _T_23720 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24388 = _T_24387 | _T_24133; // @[Mux.scala 27:72]
  wire  _T_23722 = bht_rd_addr_hashed_p1_f == 8'h64; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_100; // @[Reg.scala 27:20]
  wire [1:0] _T_24134 = _T_23722 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24389 = _T_24388 | _T_24134; // @[Mux.scala 27:72]
  wire  _T_23724 = bht_rd_addr_hashed_p1_f == 8'h65; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_101; // @[Reg.scala 27:20]
  wire [1:0] _T_24135 = _T_23724 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24390 = _T_24389 | _T_24135; // @[Mux.scala 27:72]
  wire  _T_23726 = bht_rd_addr_hashed_p1_f == 8'h66; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_102; // @[Reg.scala 27:20]
  wire [1:0] _T_24136 = _T_23726 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24391 = _T_24390 | _T_24136; // @[Mux.scala 27:72]
  wire  _T_23728 = bht_rd_addr_hashed_p1_f == 8'h67; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_103; // @[Reg.scala 27:20]
  wire [1:0] _T_24137 = _T_23728 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24392 = _T_24391 | _T_24137; // @[Mux.scala 27:72]
  wire  _T_23730 = bht_rd_addr_hashed_p1_f == 8'h68; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_104; // @[Reg.scala 27:20]
  wire [1:0] _T_24138 = _T_23730 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24393 = _T_24392 | _T_24138; // @[Mux.scala 27:72]
  wire  _T_23732 = bht_rd_addr_hashed_p1_f == 8'h69; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_105; // @[Reg.scala 27:20]
  wire [1:0] _T_24139 = _T_23732 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24394 = _T_24393 | _T_24139; // @[Mux.scala 27:72]
  wire  _T_23734 = bht_rd_addr_hashed_p1_f == 8'h6a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_106; // @[Reg.scala 27:20]
  wire [1:0] _T_24140 = _T_23734 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24395 = _T_24394 | _T_24140; // @[Mux.scala 27:72]
  wire  _T_23736 = bht_rd_addr_hashed_p1_f == 8'h6b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_107; // @[Reg.scala 27:20]
  wire [1:0] _T_24141 = _T_23736 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24396 = _T_24395 | _T_24141; // @[Mux.scala 27:72]
  wire  _T_23738 = bht_rd_addr_hashed_p1_f == 8'h6c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_108; // @[Reg.scala 27:20]
  wire [1:0] _T_24142 = _T_23738 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24397 = _T_24396 | _T_24142; // @[Mux.scala 27:72]
  wire  _T_23740 = bht_rd_addr_hashed_p1_f == 8'h6d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_109; // @[Reg.scala 27:20]
  wire [1:0] _T_24143 = _T_23740 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24398 = _T_24397 | _T_24143; // @[Mux.scala 27:72]
  wire  _T_23742 = bht_rd_addr_hashed_p1_f == 8'h6e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_110; // @[Reg.scala 27:20]
  wire [1:0] _T_24144 = _T_23742 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24399 = _T_24398 | _T_24144; // @[Mux.scala 27:72]
  wire  _T_23744 = bht_rd_addr_hashed_p1_f == 8'h6f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_111; // @[Reg.scala 27:20]
  wire [1:0] _T_24145 = _T_23744 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24400 = _T_24399 | _T_24145; // @[Mux.scala 27:72]
  wire  _T_23746 = bht_rd_addr_hashed_p1_f == 8'h70; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_112; // @[Reg.scala 27:20]
  wire [1:0] _T_24146 = _T_23746 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24401 = _T_24400 | _T_24146; // @[Mux.scala 27:72]
  wire  _T_23748 = bht_rd_addr_hashed_p1_f == 8'h71; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_113; // @[Reg.scala 27:20]
  wire [1:0] _T_24147 = _T_23748 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24402 = _T_24401 | _T_24147; // @[Mux.scala 27:72]
  wire  _T_23750 = bht_rd_addr_hashed_p1_f == 8'h72; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_114; // @[Reg.scala 27:20]
  wire [1:0] _T_24148 = _T_23750 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24403 = _T_24402 | _T_24148; // @[Mux.scala 27:72]
  wire  _T_23752 = bht_rd_addr_hashed_p1_f == 8'h73; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_115; // @[Reg.scala 27:20]
  wire [1:0] _T_24149 = _T_23752 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24404 = _T_24403 | _T_24149; // @[Mux.scala 27:72]
  wire  _T_23754 = bht_rd_addr_hashed_p1_f == 8'h74; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_116; // @[Reg.scala 27:20]
  wire [1:0] _T_24150 = _T_23754 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24405 = _T_24404 | _T_24150; // @[Mux.scala 27:72]
  wire  _T_23756 = bht_rd_addr_hashed_p1_f == 8'h75; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_117; // @[Reg.scala 27:20]
  wire [1:0] _T_24151 = _T_23756 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24406 = _T_24405 | _T_24151; // @[Mux.scala 27:72]
  wire  _T_23758 = bht_rd_addr_hashed_p1_f == 8'h76; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_118; // @[Reg.scala 27:20]
  wire [1:0] _T_24152 = _T_23758 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24407 = _T_24406 | _T_24152; // @[Mux.scala 27:72]
  wire  _T_23760 = bht_rd_addr_hashed_p1_f == 8'h77; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_119; // @[Reg.scala 27:20]
  wire [1:0] _T_24153 = _T_23760 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24408 = _T_24407 | _T_24153; // @[Mux.scala 27:72]
  wire  _T_23762 = bht_rd_addr_hashed_p1_f == 8'h78; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_120; // @[Reg.scala 27:20]
  wire [1:0] _T_24154 = _T_23762 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24409 = _T_24408 | _T_24154; // @[Mux.scala 27:72]
  wire  _T_23764 = bht_rd_addr_hashed_p1_f == 8'h79; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_121; // @[Reg.scala 27:20]
  wire [1:0] _T_24155 = _T_23764 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24410 = _T_24409 | _T_24155; // @[Mux.scala 27:72]
  wire  _T_23766 = bht_rd_addr_hashed_p1_f == 8'h7a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_122; // @[Reg.scala 27:20]
  wire [1:0] _T_24156 = _T_23766 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24411 = _T_24410 | _T_24156; // @[Mux.scala 27:72]
  wire  _T_23768 = bht_rd_addr_hashed_p1_f == 8'h7b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_123; // @[Reg.scala 27:20]
  wire [1:0] _T_24157 = _T_23768 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24412 = _T_24411 | _T_24157; // @[Mux.scala 27:72]
  wire  _T_23770 = bht_rd_addr_hashed_p1_f == 8'h7c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_124; // @[Reg.scala 27:20]
  wire [1:0] _T_24158 = _T_23770 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24413 = _T_24412 | _T_24158; // @[Mux.scala 27:72]
  wire  _T_23772 = bht_rd_addr_hashed_p1_f == 8'h7d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_125; // @[Reg.scala 27:20]
  wire [1:0] _T_24159 = _T_23772 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24414 = _T_24413 | _T_24159; // @[Mux.scala 27:72]
  wire  _T_23774 = bht_rd_addr_hashed_p1_f == 8'h7e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_126; // @[Reg.scala 27:20]
  wire [1:0] _T_24160 = _T_23774 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24415 = _T_24414 | _T_24160; // @[Mux.scala 27:72]
  wire  _T_23776 = bht_rd_addr_hashed_p1_f == 8'h7f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_127; // @[Reg.scala 27:20]
  wire [1:0] _T_24161 = _T_23776 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24416 = _T_24415 | _T_24161; // @[Mux.scala 27:72]
  wire  _T_23778 = bht_rd_addr_hashed_p1_f == 8'h80; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_128; // @[Reg.scala 27:20]
  wire [1:0] _T_24162 = _T_23778 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24417 = _T_24416 | _T_24162; // @[Mux.scala 27:72]
  wire  _T_23780 = bht_rd_addr_hashed_p1_f == 8'h81; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_129; // @[Reg.scala 27:20]
  wire [1:0] _T_24163 = _T_23780 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24418 = _T_24417 | _T_24163; // @[Mux.scala 27:72]
  wire  _T_23782 = bht_rd_addr_hashed_p1_f == 8'h82; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_130; // @[Reg.scala 27:20]
  wire [1:0] _T_24164 = _T_23782 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24419 = _T_24418 | _T_24164; // @[Mux.scala 27:72]
  wire  _T_23784 = bht_rd_addr_hashed_p1_f == 8'h83; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_131; // @[Reg.scala 27:20]
  wire [1:0] _T_24165 = _T_23784 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24420 = _T_24419 | _T_24165; // @[Mux.scala 27:72]
  wire  _T_23786 = bht_rd_addr_hashed_p1_f == 8'h84; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_132; // @[Reg.scala 27:20]
  wire [1:0] _T_24166 = _T_23786 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24421 = _T_24420 | _T_24166; // @[Mux.scala 27:72]
  wire  _T_23788 = bht_rd_addr_hashed_p1_f == 8'h85; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_133; // @[Reg.scala 27:20]
  wire [1:0] _T_24167 = _T_23788 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24422 = _T_24421 | _T_24167; // @[Mux.scala 27:72]
  wire  _T_23790 = bht_rd_addr_hashed_p1_f == 8'h86; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_134; // @[Reg.scala 27:20]
  wire [1:0] _T_24168 = _T_23790 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24423 = _T_24422 | _T_24168; // @[Mux.scala 27:72]
  wire  _T_23792 = bht_rd_addr_hashed_p1_f == 8'h87; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_135; // @[Reg.scala 27:20]
  wire [1:0] _T_24169 = _T_23792 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24424 = _T_24423 | _T_24169; // @[Mux.scala 27:72]
  wire  _T_23794 = bht_rd_addr_hashed_p1_f == 8'h88; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_136; // @[Reg.scala 27:20]
  wire [1:0] _T_24170 = _T_23794 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24425 = _T_24424 | _T_24170; // @[Mux.scala 27:72]
  wire  _T_23796 = bht_rd_addr_hashed_p1_f == 8'h89; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_137; // @[Reg.scala 27:20]
  wire [1:0] _T_24171 = _T_23796 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24426 = _T_24425 | _T_24171; // @[Mux.scala 27:72]
  wire  _T_23798 = bht_rd_addr_hashed_p1_f == 8'h8a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_138; // @[Reg.scala 27:20]
  wire [1:0] _T_24172 = _T_23798 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24427 = _T_24426 | _T_24172; // @[Mux.scala 27:72]
  wire  _T_23800 = bht_rd_addr_hashed_p1_f == 8'h8b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_139; // @[Reg.scala 27:20]
  wire [1:0] _T_24173 = _T_23800 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24428 = _T_24427 | _T_24173; // @[Mux.scala 27:72]
  wire  _T_23802 = bht_rd_addr_hashed_p1_f == 8'h8c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_140; // @[Reg.scala 27:20]
  wire [1:0] _T_24174 = _T_23802 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24429 = _T_24428 | _T_24174; // @[Mux.scala 27:72]
  wire  _T_23804 = bht_rd_addr_hashed_p1_f == 8'h8d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_141; // @[Reg.scala 27:20]
  wire [1:0] _T_24175 = _T_23804 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24430 = _T_24429 | _T_24175; // @[Mux.scala 27:72]
  wire  _T_23806 = bht_rd_addr_hashed_p1_f == 8'h8e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_142; // @[Reg.scala 27:20]
  wire [1:0] _T_24176 = _T_23806 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24431 = _T_24430 | _T_24176; // @[Mux.scala 27:72]
  wire  _T_23808 = bht_rd_addr_hashed_p1_f == 8'h8f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_143; // @[Reg.scala 27:20]
  wire [1:0] _T_24177 = _T_23808 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24432 = _T_24431 | _T_24177; // @[Mux.scala 27:72]
  wire  _T_23810 = bht_rd_addr_hashed_p1_f == 8'h90; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_144; // @[Reg.scala 27:20]
  wire [1:0] _T_24178 = _T_23810 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24433 = _T_24432 | _T_24178; // @[Mux.scala 27:72]
  wire  _T_23812 = bht_rd_addr_hashed_p1_f == 8'h91; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_145; // @[Reg.scala 27:20]
  wire [1:0] _T_24179 = _T_23812 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24434 = _T_24433 | _T_24179; // @[Mux.scala 27:72]
  wire  _T_23814 = bht_rd_addr_hashed_p1_f == 8'h92; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_146; // @[Reg.scala 27:20]
  wire [1:0] _T_24180 = _T_23814 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24435 = _T_24434 | _T_24180; // @[Mux.scala 27:72]
  wire  _T_23816 = bht_rd_addr_hashed_p1_f == 8'h93; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_147; // @[Reg.scala 27:20]
  wire [1:0] _T_24181 = _T_23816 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24436 = _T_24435 | _T_24181; // @[Mux.scala 27:72]
  wire  _T_23818 = bht_rd_addr_hashed_p1_f == 8'h94; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_148; // @[Reg.scala 27:20]
  wire [1:0] _T_24182 = _T_23818 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24437 = _T_24436 | _T_24182; // @[Mux.scala 27:72]
  wire  _T_23820 = bht_rd_addr_hashed_p1_f == 8'h95; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_149; // @[Reg.scala 27:20]
  wire [1:0] _T_24183 = _T_23820 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24438 = _T_24437 | _T_24183; // @[Mux.scala 27:72]
  wire  _T_23822 = bht_rd_addr_hashed_p1_f == 8'h96; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_150; // @[Reg.scala 27:20]
  wire [1:0] _T_24184 = _T_23822 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24439 = _T_24438 | _T_24184; // @[Mux.scala 27:72]
  wire  _T_23824 = bht_rd_addr_hashed_p1_f == 8'h97; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_151; // @[Reg.scala 27:20]
  wire [1:0] _T_24185 = _T_23824 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24440 = _T_24439 | _T_24185; // @[Mux.scala 27:72]
  wire  _T_23826 = bht_rd_addr_hashed_p1_f == 8'h98; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_152; // @[Reg.scala 27:20]
  wire [1:0] _T_24186 = _T_23826 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24441 = _T_24440 | _T_24186; // @[Mux.scala 27:72]
  wire  _T_23828 = bht_rd_addr_hashed_p1_f == 8'h99; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_153; // @[Reg.scala 27:20]
  wire [1:0] _T_24187 = _T_23828 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24442 = _T_24441 | _T_24187; // @[Mux.scala 27:72]
  wire  _T_23830 = bht_rd_addr_hashed_p1_f == 8'h9a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_154; // @[Reg.scala 27:20]
  wire [1:0] _T_24188 = _T_23830 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24443 = _T_24442 | _T_24188; // @[Mux.scala 27:72]
  wire  _T_23832 = bht_rd_addr_hashed_p1_f == 8'h9b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_155; // @[Reg.scala 27:20]
  wire [1:0] _T_24189 = _T_23832 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24444 = _T_24443 | _T_24189; // @[Mux.scala 27:72]
  wire  _T_23834 = bht_rd_addr_hashed_p1_f == 8'h9c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_156; // @[Reg.scala 27:20]
  wire [1:0] _T_24190 = _T_23834 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24445 = _T_24444 | _T_24190; // @[Mux.scala 27:72]
  wire  _T_23836 = bht_rd_addr_hashed_p1_f == 8'h9d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_157; // @[Reg.scala 27:20]
  wire [1:0] _T_24191 = _T_23836 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24446 = _T_24445 | _T_24191; // @[Mux.scala 27:72]
  wire  _T_23838 = bht_rd_addr_hashed_p1_f == 8'h9e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_158; // @[Reg.scala 27:20]
  wire [1:0] _T_24192 = _T_23838 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24447 = _T_24446 | _T_24192; // @[Mux.scala 27:72]
  wire  _T_23840 = bht_rd_addr_hashed_p1_f == 8'h9f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_159; // @[Reg.scala 27:20]
  wire [1:0] _T_24193 = _T_23840 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24448 = _T_24447 | _T_24193; // @[Mux.scala 27:72]
  wire  _T_23842 = bht_rd_addr_hashed_p1_f == 8'ha0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_160; // @[Reg.scala 27:20]
  wire [1:0] _T_24194 = _T_23842 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24449 = _T_24448 | _T_24194; // @[Mux.scala 27:72]
  wire  _T_23844 = bht_rd_addr_hashed_p1_f == 8'ha1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_161; // @[Reg.scala 27:20]
  wire [1:0] _T_24195 = _T_23844 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24450 = _T_24449 | _T_24195; // @[Mux.scala 27:72]
  wire  _T_23846 = bht_rd_addr_hashed_p1_f == 8'ha2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_162; // @[Reg.scala 27:20]
  wire [1:0] _T_24196 = _T_23846 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24451 = _T_24450 | _T_24196; // @[Mux.scala 27:72]
  wire  _T_23848 = bht_rd_addr_hashed_p1_f == 8'ha3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_163; // @[Reg.scala 27:20]
  wire [1:0] _T_24197 = _T_23848 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24452 = _T_24451 | _T_24197; // @[Mux.scala 27:72]
  wire  _T_23850 = bht_rd_addr_hashed_p1_f == 8'ha4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_164; // @[Reg.scala 27:20]
  wire [1:0] _T_24198 = _T_23850 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24453 = _T_24452 | _T_24198; // @[Mux.scala 27:72]
  wire  _T_23852 = bht_rd_addr_hashed_p1_f == 8'ha5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_165; // @[Reg.scala 27:20]
  wire [1:0] _T_24199 = _T_23852 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24454 = _T_24453 | _T_24199; // @[Mux.scala 27:72]
  wire  _T_23854 = bht_rd_addr_hashed_p1_f == 8'ha6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_166; // @[Reg.scala 27:20]
  wire [1:0] _T_24200 = _T_23854 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24455 = _T_24454 | _T_24200; // @[Mux.scala 27:72]
  wire  _T_23856 = bht_rd_addr_hashed_p1_f == 8'ha7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_167; // @[Reg.scala 27:20]
  wire [1:0] _T_24201 = _T_23856 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24456 = _T_24455 | _T_24201; // @[Mux.scala 27:72]
  wire  _T_23858 = bht_rd_addr_hashed_p1_f == 8'ha8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_168; // @[Reg.scala 27:20]
  wire [1:0] _T_24202 = _T_23858 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24457 = _T_24456 | _T_24202; // @[Mux.scala 27:72]
  wire  _T_23860 = bht_rd_addr_hashed_p1_f == 8'ha9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_169; // @[Reg.scala 27:20]
  wire [1:0] _T_24203 = _T_23860 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24458 = _T_24457 | _T_24203; // @[Mux.scala 27:72]
  wire  _T_23862 = bht_rd_addr_hashed_p1_f == 8'haa; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_170; // @[Reg.scala 27:20]
  wire [1:0] _T_24204 = _T_23862 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24459 = _T_24458 | _T_24204; // @[Mux.scala 27:72]
  wire  _T_23864 = bht_rd_addr_hashed_p1_f == 8'hab; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_171; // @[Reg.scala 27:20]
  wire [1:0] _T_24205 = _T_23864 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24460 = _T_24459 | _T_24205; // @[Mux.scala 27:72]
  wire  _T_23866 = bht_rd_addr_hashed_p1_f == 8'hac; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_172; // @[Reg.scala 27:20]
  wire [1:0] _T_24206 = _T_23866 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24461 = _T_24460 | _T_24206; // @[Mux.scala 27:72]
  wire  _T_23868 = bht_rd_addr_hashed_p1_f == 8'had; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_173; // @[Reg.scala 27:20]
  wire [1:0] _T_24207 = _T_23868 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24462 = _T_24461 | _T_24207; // @[Mux.scala 27:72]
  wire  _T_23870 = bht_rd_addr_hashed_p1_f == 8'hae; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_174; // @[Reg.scala 27:20]
  wire [1:0] _T_24208 = _T_23870 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24463 = _T_24462 | _T_24208; // @[Mux.scala 27:72]
  wire  _T_23872 = bht_rd_addr_hashed_p1_f == 8'haf; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_175; // @[Reg.scala 27:20]
  wire [1:0] _T_24209 = _T_23872 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24464 = _T_24463 | _T_24209; // @[Mux.scala 27:72]
  wire  _T_23874 = bht_rd_addr_hashed_p1_f == 8'hb0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_176; // @[Reg.scala 27:20]
  wire [1:0] _T_24210 = _T_23874 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24465 = _T_24464 | _T_24210; // @[Mux.scala 27:72]
  wire  _T_23876 = bht_rd_addr_hashed_p1_f == 8'hb1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_177; // @[Reg.scala 27:20]
  wire [1:0] _T_24211 = _T_23876 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24466 = _T_24465 | _T_24211; // @[Mux.scala 27:72]
  wire  _T_23878 = bht_rd_addr_hashed_p1_f == 8'hb2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_178; // @[Reg.scala 27:20]
  wire [1:0] _T_24212 = _T_23878 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24467 = _T_24466 | _T_24212; // @[Mux.scala 27:72]
  wire  _T_23880 = bht_rd_addr_hashed_p1_f == 8'hb3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_179; // @[Reg.scala 27:20]
  wire [1:0] _T_24213 = _T_23880 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24468 = _T_24467 | _T_24213; // @[Mux.scala 27:72]
  wire  _T_23882 = bht_rd_addr_hashed_p1_f == 8'hb4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_180; // @[Reg.scala 27:20]
  wire [1:0] _T_24214 = _T_23882 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24469 = _T_24468 | _T_24214; // @[Mux.scala 27:72]
  wire  _T_23884 = bht_rd_addr_hashed_p1_f == 8'hb5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_181; // @[Reg.scala 27:20]
  wire [1:0] _T_24215 = _T_23884 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24470 = _T_24469 | _T_24215; // @[Mux.scala 27:72]
  wire  _T_23886 = bht_rd_addr_hashed_p1_f == 8'hb6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_182; // @[Reg.scala 27:20]
  wire [1:0] _T_24216 = _T_23886 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24471 = _T_24470 | _T_24216; // @[Mux.scala 27:72]
  wire  _T_23888 = bht_rd_addr_hashed_p1_f == 8'hb7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_183; // @[Reg.scala 27:20]
  wire [1:0] _T_24217 = _T_23888 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24472 = _T_24471 | _T_24217; // @[Mux.scala 27:72]
  wire  _T_23890 = bht_rd_addr_hashed_p1_f == 8'hb8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_184; // @[Reg.scala 27:20]
  wire [1:0] _T_24218 = _T_23890 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24473 = _T_24472 | _T_24218; // @[Mux.scala 27:72]
  wire  _T_23892 = bht_rd_addr_hashed_p1_f == 8'hb9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_185; // @[Reg.scala 27:20]
  wire [1:0] _T_24219 = _T_23892 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24474 = _T_24473 | _T_24219; // @[Mux.scala 27:72]
  wire  _T_23894 = bht_rd_addr_hashed_p1_f == 8'hba; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_186; // @[Reg.scala 27:20]
  wire [1:0] _T_24220 = _T_23894 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24475 = _T_24474 | _T_24220; // @[Mux.scala 27:72]
  wire  _T_23896 = bht_rd_addr_hashed_p1_f == 8'hbb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_187; // @[Reg.scala 27:20]
  wire [1:0] _T_24221 = _T_23896 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24476 = _T_24475 | _T_24221; // @[Mux.scala 27:72]
  wire  _T_23898 = bht_rd_addr_hashed_p1_f == 8'hbc; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_188; // @[Reg.scala 27:20]
  wire [1:0] _T_24222 = _T_23898 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24477 = _T_24476 | _T_24222; // @[Mux.scala 27:72]
  wire  _T_23900 = bht_rd_addr_hashed_p1_f == 8'hbd; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_189; // @[Reg.scala 27:20]
  wire [1:0] _T_24223 = _T_23900 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24478 = _T_24477 | _T_24223; // @[Mux.scala 27:72]
  wire  _T_23902 = bht_rd_addr_hashed_p1_f == 8'hbe; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_190; // @[Reg.scala 27:20]
  wire [1:0] _T_24224 = _T_23902 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24479 = _T_24478 | _T_24224; // @[Mux.scala 27:72]
  wire  _T_23904 = bht_rd_addr_hashed_p1_f == 8'hbf; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_191; // @[Reg.scala 27:20]
  wire [1:0] _T_24225 = _T_23904 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24480 = _T_24479 | _T_24225; // @[Mux.scala 27:72]
  wire  _T_23906 = bht_rd_addr_hashed_p1_f == 8'hc0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_192; // @[Reg.scala 27:20]
  wire [1:0] _T_24226 = _T_23906 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24481 = _T_24480 | _T_24226; // @[Mux.scala 27:72]
  wire  _T_23908 = bht_rd_addr_hashed_p1_f == 8'hc1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_193; // @[Reg.scala 27:20]
  wire [1:0] _T_24227 = _T_23908 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24482 = _T_24481 | _T_24227; // @[Mux.scala 27:72]
  wire  _T_23910 = bht_rd_addr_hashed_p1_f == 8'hc2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_194; // @[Reg.scala 27:20]
  wire [1:0] _T_24228 = _T_23910 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24483 = _T_24482 | _T_24228; // @[Mux.scala 27:72]
  wire  _T_23912 = bht_rd_addr_hashed_p1_f == 8'hc3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_195; // @[Reg.scala 27:20]
  wire [1:0] _T_24229 = _T_23912 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24484 = _T_24483 | _T_24229; // @[Mux.scala 27:72]
  wire  _T_23914 = bht_rd_addr_hashed_p1_f == 8'hc4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_196; // @[Reg.scala 27:20]
  wire [1:0] _T_24230 = _T_23914 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24485 = _T_24484 | _T_24230; // @[Mux.scala 27:72]
  wire  _T_23916 = bht_rd_addr_hashed_p1_f == 8'hc5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_197; // @[Reg.scala 27:20]
  wire [1:0] _T_24231 = _T_23916 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24486 = _T_24485 | _T_24231; // @[Mux.scala 27:72]
  wire  _T_23918 = bht_rd_addr_hashed_p1_f == 8'hc6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_198; // @[Reg.scala 27:20]
  wire [1:0] _T_24232 = _T_23918 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24487 = _T_24486 | _T_24232; // @[Mux.scala 27:72]
  wire  _T_23920 = bht_rd_addr_hashed_p1_f == 8'hc7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_199; // @[Reg.scala 27:20]
  wire [1:0] _T_24233 = _T_23920 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24488 = _T_24487 | _T_24233; // @[Mux.scala 27:72]
  wire  _T_23922 = bht_rd_addr_hashed_p1_f == 8'hc8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_200; // @[Reg.scala 27:20]
  wire [1:0] _T_24234 = _T_23922 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24489 = _T_24488 | _T_24234; // @[Mux.scala 27:72]
  wire  _T_23924 = bht_rd_addr_hashed_p1_f == 8'hc9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_201; // @[Reg.scala 27:20]
  wire [1:0] _T_24235 = _T_23924 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24490 = _T_24489 | _T_24235; // @[Mux.scala 27:72]
  wire  _T_23926 = bht_rd_addr_hashed_p1_f == 8'hca; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_202; // @[Reg.scala 27:20]
  wire [1:0] _T_24236 = _T_23926 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24491 = _T_24490 | _T_24236; // @[Mux.scala 27:72]
  wire  _T_23928 = bht_rd_addr_hashed_p1_f == 8'hcb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_203; // @[Reg.scala 27:20]
  wire [1:0] _T_24237 = _T_23928 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24492 = _T_24491 | _T_24237; // @[Mux.scala 27:72]
  wire  _T_23930 = bht_rd_addr_hashed_p1_f == 8'hcc; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_204; // @[Reg.scala 27:20]
  wire [1:0] _T_24238 = _T_23930 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24493 = _T_24492 | _T_24238; // @[Mux.scala 27:72]
  wire  _T_23932 = bht_rd_addr_hashed_p1_f == 8'hcd; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_205; // @[Reg.scala 27:20]
  wire [1:0] _T_24239 = _T_23932 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24494 = _T_24493 | _T_24239; // @[Mux.scala 27:72]
  wire  _T_23934 = bht_rd_addr_hashed_p1_f == 8'hce; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_206; // @[Reg.scala 27:20]
  wire [1:0] _T_24240 = _T_23934 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24495 = _T_24494 | _T_24240; // @[Mux.scala 27:72]
  wire  _T_23936 = bht_rd_addr_hashed_p1_f == 8'hcf; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_207; // @[Reg.scala 27:20]
  wire [1:0] _T_24241 = _T_23936 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24496 = _T_24495 | _T_24241; // @[Mux.scala 27:72]
  wire  _T_23938 = bht_rd_addr_hashed_p1_f == 8'hd0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_208; // @[Reg.scala 27:20]
  wire [1:0] _T_24242 = _T_23938 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24497 = _T_24496 | _T_24242; // @[Mux.scala 27:72]
  wire  _T_23940 = bht_rd_addr_hashed_p1_f == 8'hd1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_209; // @[Reg.scala 27:20]
  wire [1:0] _T_24243 = _T_23940 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24498 = _T_24497 | _T_24243; // @[Mux.scala 27:72]
  wire  _T_23942 = bht_rd_addr_hashed_p1_f == 8'hd2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_210; // @[Reg.scala 27:20]
  wire [1:0] _T_24244 = _T_23942 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24499 = _T_24498 | _T_24244; // @[Mux.scala 27:72]
  wire  _T_23944 = bht_rd_addr_hashed_p1_f == 8'hd3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_211; // @[Reg.scala 27:20]
  wire [1:0] _T_24245 = _T_23944 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24500 = _T_24499 | _T_24245; // @[Mux.scala 27:72]
  wire  _T_23946 = bht_rd_addr_hashed_p1_f == 8'hd4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_212; // @[Reg.scala 27:20]
  wire [1:0] _T_24246 = _T_23946 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24501 = _T_24500 | _T_24246; // @[Mux.scala 27:72]
  wire  _T_23948 = bht_rd_addr_hashed_p1_f == 8'hd5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_213; // @[Reg.scala 27:20]
  wire [1:0] _T_24247 = _T_23948 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24502 = _T_24501 | _T_24247; // @[Mux.scala 27:72]
  wire  _T_23950 = bht_rd_addr_hashed_p1_f == 8'hd6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_214; // @[Reg.scala 27:20]
  wire [1:0] _T_24248 = _T_23950 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24503 = _T_24502 | _T_24248; // @[Mux.scala 27:72]
  wire  _T_23952 = bht_rd_addr_hashed_p1_f == 8'hd7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_215; // @[Reg.scala 27:20]
  wire [1:0] _T_24249 = _T_23952 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24504 = _T_24503 | _T_24249; // @[Mux.scala 27:72]
  wire  _T_23954 = bht_rd_addr_hashed_p1_f == 8'hd8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_216; // @[Reg.scala 27:20]
  wire [1:0] _T_24250 = _T_23954 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24505 = _T_24504 | _T_24250; // @[Mux.scala 27:72]
  wire  _T_23956 = bht_rd_addr_hashed_p1_f == 8'hd9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_217; // @[Reg.scala 27:20]
  wire [1:0] _T_24251 = _T_23956 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24506 = _T_24505 | _T_24251; // @[Mux.scala 27:72]
  wire  _T_23958 = bht_rd_addr_hashed_p1_f == 8'hda; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_218; // @[Reg.scala 27:20]
  wire [1:0] _T_24252 = _T_23958 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24507 = _T_24506 | _T_24252; // @[Mux.scala 27:72]
  wire  _T_23960 = bht_rd_addr_hashed_p1_f == 8'hdb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_219; // @[Reg.scala 27:20]
  wire [1:0] _T_24253 = _T_23960 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24508 = _T_24507 | _T_24253; // @[Mux.scala 27:72]
  wire  _T_23962 = bht_rd_addr_hashed_p1_f == 8'hdc; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_220; // @[Reg.scala 27:20]
  wire [1:0] _T_24254 = _T_23962 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24509 = _T_24508 | _T_24254; // @[Mux.scala 27:72]
  wire  _T_23964 = bht_rd_addr_hashed_p1_f == 8'hdd; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_221; // @[Reg.scala 27:20]
  wire [1:0] _T_24255 = _T_23964 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24510 = _T_24509 | _T_24255; // @[Mux.scala 27:72]
  wire  _T_23966 = bht_rd_addr_hashed_p1_f == 8'hde; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_222; // @[Reg.scala 27:20]
  wire [1:0] _T_24256 = _T_23966 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24511 = _T_24510 | _T_24256; // @[Mux.scala 27:72]
  wire  _T_23968 = bht_rd_addr_hashed_p1_f == 8'hdf; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_223; // @[Reg.scala 27:20]
  wire [1:0] _T_24257 = _T_23968 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24512 = _T_24511 | _T_24257; // @[Mux.scala 27:72]
  wire  _T_23970 = bht_rd_addr_hashed_p1_f == 8'he0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_224; // @[Reg.scala 27:20]
  wire [1:0] _T_24258 = _T_23970 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24513 = _T_24512 | _T_24258; // @[Mux.scala 27:72]
  wire  _T_23972 = bht_rd_addr_hashed_p1_f == 8'he1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_225; // @[Reg.scala 27:20]
  wire [1:0] _T_24259 = _T_23972 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24514 = _T_24513 | _T_24259; // @[Mux.scala 27:72]
  wire  _T_23974 = bht_rd_addr_hashed_p1_f == 8'he2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_226; // @[Reg.scala 27:20]
  wire [1:0] _T_24260 = _T_23974 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24515 = _T_24514 | _T_24260; // @[Mux.scala 27:72]
  wire  _T_23976 = bht_rd_addr_hashed_p1_f == 8'he3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_227; // @[Reg.scala 27:20]
  wire [1:0] _T_24261 = _T_23976 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24516 = _T_24515 | _T_24261; // @[Mux.scala 27:72]
  wire  _T_23978 = bht_rd_addr_hashed_p1_f == 8'he4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_228; // @[Reg.scala 27:20]
  wire [1:0] _T_24262 = _T_23978 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24517 = _T_24516 | _T_24262; // @[Mux.scala 27:72]
  wire  _T_23980 = bht_rd_addr_hashed_p1_f == 8'he5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_229; // @[Reg.scala 27:20]
  wire [1:0] _T_24263 = _T_23980 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24518 = _T_24517 | _T_24263; // @[Mux.scala 27:72]
  wire  _T_23982 = bht_rd_addr_hashed_p1_f == 8'he6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_230; // @[Reg.scala 27:20]
  wire [1:0] _T_24264 = _T_23982 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24519 = _T_24518 | _T_24264; // @[Mux.scala 27:72]
  wire  _T_23984 = bht_rd_addr_hashed_p1_f == 8'he7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_231; // @[Reg.scala 27:20]
  wire [1:0] _T_24265 = _T_23984 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24520 = _T_24519 | _T_24265; // @[Mux.scala 27:72]
  wire  _T_23986 = bht_rd_addr_hashed_p1_f == 8'he8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_232; // @[Reg.scala 27:20]
  wire [1:0] _T_24266 = _T_23986 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24521 = _T_24520 | _T_24266; // @[Mux.scala 27:72]
  wire  _T_23988 = bht_rd_addr_hashed_p1_f == 8'he9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_233; // @[Reg.scala 27:20]
  wire [1:0] _T_24267 = _T_23988 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24522 = _T_24521 | _T_24267; // @[Mux.scala 27:72]
  wire  _T_23990 = bht_rd_addr_hashed_p1_f == 8'hea; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_234; // @[Reg.scala 27:20]
  wire [1:0] _T_24268 = _T_23990 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24523 = _T_24522 | _T_24268; // @[Mux.scala 27:72]
  wire  _T_23992 = bht_rd_addr_hashed_p1_f == 8'heb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_235; // @[Reg.scala 27:20]
  wire [1:0] _T_24269 = _T_23992 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24524 = _T_24523 | _T_24269; // @[Mux.scala 27:72]
  wire  _T_23994 = bht_rd_addr_hashed_p1_f == 8'hec; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_236; // @[Reg.scala 27:20]
  wire [1:0] _T_24270 = _T_23994 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24525 = _T_24524 | _T_24270; // @[Mux.scala 27:72]
  wire  _T_23996 = bht_rd_addr_hashed_p1_f == 8'hed; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_237; // @[Reg.scala 27:20]
  wire [1:0] _T_24271 = _T_23996 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24526 = _T_24525 | _T_24271; // @[Mux.scala 27:72]
  wire  _T_23998 = bht_rd_addr_hashed_p1_f == 8'hee; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_238; // @[Reg.scala 27:20]
  wire [1:0] _T_24272 = _T_23998 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24527 = _T_24526 | _T_24272; // @[Mux.scala 27:72]
  wire  _T_24000 = bht_rd_addr_hashed_p1_f == 8'hef; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_239; // @[Reg.scala 27:20]
  wire [1:0] _T_24273 = _T_24000 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24528 = _T_24527 | _T_24273; // @[Mux.scala 27:72]
  wire  _T_24002 = bht_rd_addr_hashed_p1_f == 8'hf0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_240; // @[Reg.scala 27:20]
  wire [1:0] _T_24274 = _T_24002 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24529 = _T_24528 | _T_24274; // @[Mux.scala 27:72]
  wire  _T_24004 = bht_rd_addr_hashed_p1_f == 8'hf1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_241; // @[Reg.scala 27:20]
  wire [1:0] _T_24275 = _T_24004 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24530 = _T_24529 | _T_24275; // @[Mux.scala 27:72]
  wire  _T_24006 = bht_rd_addr_hashed_p1_f == 8'hf2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_242; // @[Reg.scala 27:20]
  wire [1:0] _T_24276 = _T_24006 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24531 = _T_24530 | _T_24276; // @[Mux.scala 27:72]
  wire  _T_24008 = bht_rd_addr_hashed_p1_f == 8'hf3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_243; // @[Reg.scala 27:20]
  wire [1:0] _T_24277 = _T_24008 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24532 = _T_24531 | _T_24277; // @[Mux.scala 27:72]
  wire  _T_24010 = bht_rd_addr_hashed_p1_f == 8'hf4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_244; // @[Reg.scala 27:20]
  wire [1:0] _T_24278 = _T_24010 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24533 = _T_24532 | _T_24278; // @[Mux.scala 27:72]
  wire  _T_24012 = bht_rd_addr_hashed_p1_f == 8'hf5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_245; // @[Reg.scala 27:20]
  wire [1:0] _T_24279 = _T_24012 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24534 = _T_24533 | _T_24279; // @[Mux.scala 27:72]
  wire  _T_24014 = bht_rd_addr_hashed_p1_f == 8'hf6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_246; // @[Reg.scala 27:20]
  wire [1:0] _T_24280 = _T_24014 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24535 = _T_24534 | _T_24280; // @[Mux.scala 27:72]
  wire  _T_24016 = bht_rd_addr_hashed_p1_f == 8'hf7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_247; // @[Reg.scala 27:20]
  wire [1:0] _T_24281 = _T_24016 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24536 = _T_24535 | _T_24281; // @[Mux.scala 27:72]
  wire  _T_24018 = bht_rd_addr_hashed_p1_f == 8'hf8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_248; // @[Reg.scala 27:20]
  wire [1:0] _T_24282 = _T_24018 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24537 = _T_24536 | _T_24282; // @[Mux.scala 27:72]
  wire  _T_24020 = bht_rd_addr_hashed_p1_f == 8'hf9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_249; // @[Reg.scala 27:20]
  wire [1:0] _T_24283 = _T_24020 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24538 = _T_24537 | _T_24283; // @[Mux.scala 27:72]
  wire  _T_24022 = bht_rd_addr_hashed_p1_f == 8'hfa; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_250; // @[Reg.scala 27:20]
  wire [1:0] _T_24284 = _T_24022 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24539 = _T_24538 | _T_24284; // @[Mux.scala 27:72]
  wire  _T_24024 = bht_rd_addr_hashed_p1_f == 8'hfb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_251; // @[Reg.scala 27:20]
  wire [1:0] _T_24285 = _T_24024 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24540 = _T_24539 | _T_24285; // @[Mux.scala 27:72]
  wire  _T_24026 = bht_rd_addr_hashed_p1_f == 8'hfc; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_252; // @[Reg.scala 27:20]
  wire [1:0] _T_24286 = _T_24026 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24541 = _T_24540 | _T_24286; // @[Mux.scala 27:72]
  wire  _T_24028 = bht_rd_addr_hashed_p1_f == 8'hfd; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_253; // @[Reg.scala 27:20]
  wire [1:0] _T_24287 = _T_24028 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24542 = _T_24541 | _T_24287; // @[Mux.scala 27:72]
  wire  _T_24030 = bht_rd_addr_hashed_p1_f == 8'hfe; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_254; // @[Reg.scala 27:20]
  wire [1:0] _T_24288 = _T_24030 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24543 = _T_24542 | _T_24288; // @[Mux.scala 27:72]
  wire  _T_24032 = bht_rd_addr_hashed_p1_f == 8'hff; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_255; // @[Reg.scala 27:20]
  wire [1:0] _T_24289 = _T_24032 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_p1_f = _T_24543 | _T_24289; // @[Mux.scala 27:72]
  wire [1:0] _T_280 = io_ifc_fetch_addr_f[0] ? bht_bank0_rd_data_p1_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank1_rd_data_f = _T_279 | _T_280; // @[Mux.scala 27:72]
  wire  _T_284 = bht_force_taken_f[1] | bht_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 298:42]
  wire [1:0] wayhit_f = _T_97 | _T_107; // @[ifu_bp_ctl.scala 172:41]
  wire [1:0] _T_636 = _T_162 ? wayhit_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] wayhit_p1_f = _T_117 | _T_127; // @[ifu_bp_ctl.scala 174:47]
  wire [1:0] _T_635 = {wayhit_p1_f[0],wayhit_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_637 = io_ifc_fetch_addr_f[0] ? _T_635 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_638 = _T_636 | _T_637; // @[Mux.scala 27:72]
  wire  eoc_near = &io_ifc_fetch_addr_f[4:2]; // @[ifu_bp_ctl.scala 258:64]
  wire  _T_238 = ~eoc_near; // @[ifu_bp_ctl.scala 260:15]
  wire [1:0] _T_240 = ~io_ifc_fetch_addr_f[1:0]; // @[ifu_bp_ctl.scala 260:28]
  wire  _T_241 = |_T_240; // @[ifu_bp_ctl.scala 260:58]
  wire  eoc_mask = _T_238 | _T_241; // @[ifu_bp_ctl.scala 260:25]
  wire [1:0] _T_640 = {eoc_mask,1'h1}; // @[Cat.scala 29:58]
  wire [1:0] bht_valid_f = _T_638 & _T_640; // @[ifu_bp_ctl.scala 431:71]
  wire  _T_286 = _T_284 & bht_valid_f[1]; // @[ifu_bp_ctl.scala 298:69]
  wire [1:0] _T_21986 = _T_22498 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21987 = _T_22500 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22242 = _T_21986 | _T_21987; // @[Mux.scala 27:72]
  wire [1:0] _T_21988 = _T_22502 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22243 = _T_22242 | _T_21988; // @[Mux.scala 27:72]
  wire [1:0] _T_21989 = _T_22504 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22244 = _T_22243 | _T_21989; // @[Mux.scala 27:72]
  wire [1:0] _T_21990 = _T_22506 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22245 = _T_22244 | _T_21990; // @[Mux.scala 27:72]
  wire [1:0] _T_21991 = _T_22508 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22246 = _T_22245 | _T_21991; // @[Mux.scala 27:72]
  wire [1:0] _T_21992 = _T_22510 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22247 = _T_22246 | _T_21992; // @[Mux.scala 27:72]
  wire [1:0] _T_21993 = _T_22512 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22248 = _T_22247 | _T_21993; // @[Mux.scala 27:72]
  wire [1:0] _T_21994 = _T_22514 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22249 = _T_22248 | _T_21994; // @[Mux.scala 27:72]
  wire [1:0] _T_21995 = _T_22516 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22250 = _T_22249 | _T_21995; // @[Mux.scala 27:72]
  wire [1:0] _T_21996 = _T_22518 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22251 = _T_22250 | _T_21996; // @[Mux.scala 27:72]
  wire [1:0] _T_21997 = _T_22520 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22252 = _T_22251 | _T_21997; // @[Mux.scala 27:72]
  wire [1:0] _T_21998 = _T_22522 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22253 = _T_22252 | _T_21998; // @[Mux.scala 27:72]
  wire [1:0] _T_21999 = _T_22524 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22254 = _T_22253 | _T_21999; // @[Mux.scala 27:72]
  wire [1:0] _T_22000 = _T_22526 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22255 = _T_22254 | _T_22000; // @[Mux.scala 27:72]
  wire [1:0] _T_22001 = _T_22528 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22256 = _T_22255 | _T_22001; // @[Mux.scala 27:72]
  wire [1:0] _T_22002 = _T_22530 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22257 = _T_22256 | _T_22002; // @[Mux.scala 27:72]
  wire [1:0] _T_22003 = _T_22532 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22258 = _T_22257 | _T_22003; // @[Mux.scala 27:72]
  wire [1:0] _T_22004 = _T_22534 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22259 = _T_22258 | _T_22004; // @[Mux.scala 27:72]
  wire [1:0] _T_22005 = _T_22536 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22260 = _T_22259 | _T_22005; // @[Mux.scala 27:72]
  wire [1:0] _T_22006 = _T_22538 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22261 = _T_22260 | _T_22006; // @[Mux.scala 27:72]
  wire [1:0] _T_22007 = _T_22540 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22262 = _T_22261 | _T_22007; // @[Mux.scala 27:72]
  wire [1:0] _T_22008 = _T_22542 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22263 = _T_22262 | _T_22008; // @[Mux.scala 27:72]
  wire [1:0] _T_22009 = _T_22544 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22264 = _T_22263 | _T_22009; // @[Mux.scala 27:72]
  wire [1:0] _T_22010 = _T_22546 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22265 = _T_22264 | _T_22010; // @[Mux.scala 27:72]
  wire [1:0] _T_22011 = _T_22548 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22266 = _T_22265 | _T_22011; // @[Mux.scala 27:72]
  wire [1:0] _T_22012 = _T_22550 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22267 = _T_22266 | _T_22012; // @[Mux.scala 27:72]
  wire [1:0] _T_22013 = _T_22552 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22268 = _T_22267 | _T_22013; // @[Mux.scala 27:72]
  wire [1:0] _T_22014 = _T_22554 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22269 = _T_22268 | _T_22014; // @[Mux.scala 27:72]
  wire [1:0] _T_22015 = _T_22556 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22270 = _T_22269 | _T_22015; // @[Mux.scala 27:72]
  wire [1:0] _T_22016 = _T_22558 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22271 = _T_22270 | _T_22016; // @[Mux.scala 27:72]
  wire [1:0] _T_22017 = _T_22560 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22272 = _T_22271 | _T_22017; // @[Mux.scala 27:72]
  wire [1:0] _T_22018 = _T_22562 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22273 = _T_22272 | _T_22018; // @[Mux.scala 27:72]
  wire [1:0] _T_22019 = _T_22564 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22274 = _T_22273 | _T_22019; // @[Mux.scala 27:72]
  wire [1:0] _T_22020 = _T_22566 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22275 = _T_22274 | _T_22020; // @[Mux.scala 27:72]
  wire [1:0] _T_22021 = _T_22568 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22276 = _T_22275 | _T_22021; // @[Mux.scala 27:72]
  wire [1:0] _T_22022 = _T_22570 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22277 = _T_22276 | _T_22022; // @[Mux.scala 27:72]
  wire [1:0] _T_22023 = _T_22572 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22278 = _T_22277 | _T_22023; // @[Mux.scala 27:72]
  wire [1:0] _T_22024 = _T_22574 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22279 = _T_22278 | _T_22024; // @[Mux.scala 27:72]
  wire [1:0] _T_22025 = _T_22576 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22280 = _T_22279 | _T_22025; // @[Mux.scala 27:72]
  wire [1:0] _T_22026 = _T_22578 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22281 = _T_22280 | _T_22026; // @[Mux.scala 27:72]
  wire [1:0] _T_22027 = _T_22580 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22282 = _T_22281 | _T_22027; // @[Mux.scala 27:72]
  wire [1:0] _T_22028 = _T_22582 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22283 = _T_22282 | _T_22028; // @[Mux.scala 27:72]
  wire [1:0] _T_22029 = _T_22584 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22284 = _T_22283 | _T_22029; // @[Mux.scala 27:72]
  wire [1:0] _T_22030 = _T_22586 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22285 = _T_22284 | _T_22030; // @[Mux.scala 27:72]
  wire [1:0] _T_22031 = _T_22588 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22286 = _T_22285 | _T_22031; // @[Mux.scala 27:72]
  wire [1:0] _T_22032 = _T_22590 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22287 = _T_22286 | _T_22032; // @[Mux.scala 27:72]
  wire [1:0] _T_22033 = _T_22592 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22288 = _T_22287 | _T_22033; // @[Mux.scala 27:72]
  wire [1:0] _T_22034 = _T_22594 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22289 = _T_22288 | _T_22034; // @[Mux.scala 27:72]
  wire [1:0] _T_22035 = _T_22596 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22290 = _T_22289 | _T_22035; // @[Mux.scala 27:72]
  wire [1:0] _T_22036 = _T_22598 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22291 = _T_22290 | _T_22036; // @[Mux.scala 27:72]
  wire [1:0] _T_22037 = _T_22600 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22292 = _T_22291 | _T_22037; // @[Mux.scala 27:72]
  wire [1:0] _T_22038 = _T_22602 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22293 = _T_22292 | _T_22038; // @[Mux.scala 27:72]
  wire [1:0] _T_22039 = _T_22604 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22294 = _T_22293 | _T_22039; // @[Mux.scala 27:72]
  wire [1:0] _T_22040 = _T_22606 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22295 = _T_22294 | _T_22040; // @[Mux.scala 27:72]
  wire [1:0] _T_22041 = _T_22608 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22296 = _T_22295 | _T_22041; // @[Mux.scala 27:72]
  wire [1:0] _T_22042 = _T_22610 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22297 = _T_22296 | _T_22042; // @[Mux.scala 27:72]
  wire [1:0] _T_22043 = _T_22612 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22298 = _T_22297 | _T_22043; // @[Mux.scala 27:72]
  wire [1:0] _T_22044 = _T_22614 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22299 = _T_22298 | _T_22044; // @[Mux.scala 27:72]
  wire [1:0] _T_22045 = _T_22616 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22300 = _T_22299 | _T_22045; // @[Mux.scala 27:72]
  wire [1:0] _T_22046 = _T_22618 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22301 = _T_22300 | _T_22046; // @[Mux.scala 27:72]
  wire [1:0] _T_22047 = _T_22620 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22302 = _T_22301 | _T_22047; // @[Mux.scala 27:72]
  wire [1:0] _T_22048 = _T_22622 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22303 = _T_22302 | _T_22048; // @[Mux.scala 27:72]
  wire [1:0] _T_22049 = _T_22624 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22304 = _T_22303 | _T_22049; // @[Mux.scala 27:72]
  wire [1:0] _T_22050 = _T_22626 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22305 = _T_22304 | _T_22050; // @[Mux.scala 27:72]
  wire [1:0] _T_22051 = _T_22628 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22306 = _T_22305 | _T_22051; // @[Mux.scala 27:72]
  wire [1:0] _T_22052 = _T_22630 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22307 = _T_22306 | _T_22052; // @[Mux.scala 27:72]
  wire [1:0] _T_22053 = _T_22632 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22308 = _T_22307 | _T_22053; // @[Mux.scala 27:72]
  wire [1:0] _T_22054 = _T_22634 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22309 = _T_22308 | _T_22054; // @[Mux.scala 27:72]
  wire [1:0] _T_22055 = _T_22636 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22310 = _T_22309 | _T_22055; // @[Mux.scala 27:72]
  wire [1:0] _T_22056 = _T_22638 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22311 = _T_22310 | _T_22056; // @[Mux.scala 27:72]
  wire [1:0] _T_22057 = _T_22640 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22312 = _T_22311 | _T_22057; // @[Mux.scala 27:72]
  wire [1:0] _T_22058 = _T_22642 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22313 = _T_22312 | _T_22058; // @[Mux.scala 27:72]
  wire [1:0] _T_22059 = _T_22644 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22314 = _T_22313 | _T_22059; // @[Mux.scala 27:72]
  wire [1:0] _T_22060 = _T_22646 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22315 = _T_22314 | _T_22060; // @[Mux.scala 27:72]
  wire [1:0] _T_22061 = _T_22648 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22316 = _T_22315 | _T_22061; // @[Mux.scala 27:72]
  wire [1:0] _T_22062 = _T_22650 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22317 = _T_22316 | _T_22062; // @[Mux.scala 27:72]
  wire [1:0] _T_22063 = _T_22652 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22318 = _T_22317 | _T_22063; // @[Mux.scala 27:72]
  wire [1:0] _T_22064 = _T_22654 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22319 = _T_22318 | _T_22064; // @[Mux.scala 27:72]
  wire [1:0] _T_22065 = _T_22656 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22320 = _T_22319 | _T_22065; // @[Mux.scala 27:72]
  wire [1:0] _T_22066 = _T_22658 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22321 = _T_22320 | _T_22066; // @[Mux.scala 27:72]
  wire [1:0] _T_22067 = _T_22660 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22322 = _T_22321 | _T_22067; // @[Mux.scala 27:72]
  wire [1:0] _T_22068 = _T_22662 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22323 = _T_22322 | _T_22068; // @[Mux.scala 27:72]
  wire [1:0] _T_22069 = _T_22664 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22324 = _T_22323 | _T_22069; // @[Mux.scala 27:72]
  wire [1:0] _T_22070 = _T_22666 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22325 = _T_22324 | _T_22070; // @[Mux.scala 27:72]
  wire [1:0] _T_22071 = _T_22668 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22326 = _T_22325 | _T_22071; // @[Mux.scala 27:72]
  wire [1:0] _T_22072 = _T_22670 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22327 = _T_22326 | _T_22072; // @[Mux.scala 27:72]
  wire [1:0] _T_22073 = _T_22672 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22328 = _T_22327 | _T_22073; // @[Mux.scala 27:72]
  wire [1:0] _T_22074 = _T_22674 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22329 = _T_22328 | _T_22074; // @[Mux.scala 27:72]
  wire [1:0] _T_22075 = _T_22676 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22330 = _T_22329 | _T_22075; // @[Mux.scala 27:72]
  wire [1:0] _T_22076 = _T_22678 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22331 = _T_22330 | _T_22076; // @[Mux.scala 27:72]
  wire [1:0] _T_22077 = _T_22680 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22332 = _T_22331 | _T_22077; // @[Mux.scala 27:72]
  wire [1:0] _T_22078 = _T_22682 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22333 = _T_22332 | _T_22078; // @[Mux.scala 27:72]
  wire [1:0] _T_22079 = _T_22684 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22334 = _T_22333 | _T_22079; // @[Mux.scala 27:72]
  wire [1:0] _T_22080 = _T_22686 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22335 = _T_22334 | _T_22080; // @[Mux.scala 27:72]
  wire [1:0] _T_22081 = _T_22688 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22336 = _T_22335 | _T_22081; // @[Mux.scala 27:72]
  wire [1:0] _T_22082 = _T_22690 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22337 = _T_22336 | _T_22082; // @[Mux.scala 27:72]
  wire [1:0] _T_22083 = _T_22692 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22338 = _T_22337 | _T_22083; // @[Mux.scala 27:72]
  wire [1:0] _T_22084 = _T_22694 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22339 = _T_22338 | _T_22084; // @[Mux.scala 27:72]
  wire [1:0] _T_22085 = _T_22696 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22340 = _T_22339 | _T_22085; // @[Mux.scala 27:72]
  wire [1:0] _T_22086 = _T_22698 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22341 = _T_22340 | _T_22086; // @[Mux.scala 27:72]
  wire [1:0] _T_22087 = _T_22700 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22342 = _T_22341 | _T_22087; // @[Mux.scala 27:72]
  wire [1:0] _T_22088 = _T_22702 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22343 = _T_22342 | _T_22088; // @[Mux.scala 27:72]
  wire [1:0] _T_22089 = _T_22704 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22344 = _T_22343 | _T_22089; // @[Mux.scala 27:72]
  wire [1:0] _T_22090 = _T_22706 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22345 = _T_22344 | _T_22090; // @[Mux.scala 27:72]
  wire [1:0] _T_22091 = _T_22708 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22346 = _T_22345 | _T_22091; // @[Mux.scala 27:72]
  wire [1:0] _T_22092 = _T_22710 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22347 = _T_22346 | _T_22092; // @[Mux.scala 27:72]
  wire [1:0] _T_22093 = _T_22712 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22348 = _T_22347 | _T_22093; // @[Mux.scala 27:72]
  wire [1:0] _T_22094 = _T_22714 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22349 = _T_22348 | _T_22094; // @[Mux.scala 27:72]
  wire [1:0] _T_22095 = _T_22716 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22350 = _T_22349 | _T_22095; // @[Mux.scala 27:72]
  wire [1:0] _T_22096 = _T_22718 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22351 = _T_22350 | _T_22096; // @[Mux.scala 27:72]
  wire [1:0] _T_22097 = _T_22720 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22352 = _T_22351 | _T_22097; // @[Mux.scala 27:72]
  wire [1:0] _T_22098 = _T_22722 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22353 = _T_22352 | _T_22098; // @[Mux.scala 27:72]
  wire [1:0] _T_22099 = _T_22724 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22354 = _T_22353 | _T_22099; // @[Mux.scala 27:72]
  wire [1:0] _T_22100 = _T_22726 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22355 = _T_22354 | _T_22100; // @[Mux.scala 27:72]
  wire [1:0] _T_22101 = _T_22728 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22356 = _T_22355 | _T_22101; // @[Mux.scala 27:72]
  wire [1:0] _T_22102 = _T_22730 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22357 = _T_22356 | _T_22102; // @[Mux.scala 27:72]
  wire [1:0] _T_22103 = _T_22732 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22358 = _T_22357 | _T_22103; // @[Mux.scala 27:72]
  wire [1:0] _T_22104 = _T_22734 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22359 = _T_22358 | _T_22104; // @[Mux.scala 27:72]
  wire [1:0] _T_22105 = _T_22736 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22360 = _T_22359 | _T_22105; // @[Mux.scala 27:72]
  wire [1:0] _T_22106 = _T_22738 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22361 = _T_22360 | _T_22106; // @[Mux.scala 27:72]
  wire [1:0] _T_22107 = _T_22740 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22362 = _T_22361 | _T_22107; // @[Mux.scala 27:72]
  wire [1:0] _T_22108 = _T_22742 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22363 = _T_22362 | _T_22108; // @[Mux.scala 27:72]
  wire [1:0] _T_22109 = _T_22744 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22364 = _T_22363 | _T_22109; // @[Mux.scala 27:72]
  wire [1:0] _T_22110 = _T_22746 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22365 = _T_22364 | _T_22110; // @[Mux.scala 27:72]
  wire [1:0] _T_22111 = _T_22748 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22366 = _T_22365 | _T_22111; // @[Mux.scala 27:72]
  wire [1:0] _T_22112 = _T_22750 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22367 = _T_22366 | _T_22112; // @[Mux.scala 27:72]
  wire [1:0] _T_22113 = _T_22752 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22368 = _T_22367 | _T_22113; // @[Mux.scala 27:72]
  wire [1:0] _T_22114 = _T_22754 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22369 = _T_22368 | _T_22114; // @[Mux.scala 27:72]
  wire [1:0] _T_22115 = _T_22756 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22370 = _T_22369 | _T_22115; // @[Mux.scala 27:72]
  wire [1:0] _T_22116 = _T_22758 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22371 = _T_22370 | _T_22116; // @[Mux.scala 27:72]
  wire [1:0] _T_22117 = _T_22760 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22372 = _T_22371 | _T_22117; // @[Mux.scala 27:72]
  wire [1:0] _T_22118 = _T_22762 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22373 = _T_22372 | _T_22118; // @[Mux.scala 27:72]
  wire [1:0] _T_22119 = _T_22764 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22374 = _T_22373 | _T_22119; // @[Mux.scala 27:72]
  wire [1:0] _T_22120 = _T_22766 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22375 = _T_22374 | _T_22120; // @[Mux.scala 27:72]
  wire [1:0] _T_22121 = _T_22768 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22376 = _T_22375 | _T_22121; // @[Mux.scala 27:72]
  wire [1:0] _T_22122 = _T_22770 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22377 = _T_22376 | _T_22122; // @[Mux.scala 27:72]
  wire [1:0] _T_22123 = _T_22772 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22378 = _T_22377 | _T_22123; // @[Mux.scala 27:72]
  wire [1:0] _T_22124 = _T_22774 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22379 = _T_22378 | _T_22124; // @[Mux.scala 27:72]
  wire [1:0] _T_22125 = _T_22776 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22380 = _T_22379 | _T_22125; // @[Mux.scala 27:72]
  wire [1:0] _T_22126 = _T_22778 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22381 = _T_22380 | _T_22126; // @[Mux.scala 27:72]
  wire [1:0] _T_22127 = _T_22780 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22382 = _T_22381 | _T_22127; // @[Mux.scala 27:72]
  wire [1:0] _T_22128 = _T_22782 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22383 = _T_22382 | _T_22128; // @[Mux.scala 27:72]
  wire [1:0] _T_22129 = _T_22784 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22384 = _T_22383 | _T_22129; // @[Mux.scala 27:72]
  wire [1:0] _T_22130 = _T_22786 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22385 = _T_22384 | _T_22130; // @[Mux.scala 27:72]
  wire [1:0] _T_22131 = _T_22788 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22386 = _T_22385 | _T_22131; // @[Mux.scala 27:72]
  wire [1:0] _T_22132 = _T_22790 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22387 = _T_22386 | _T_22132; // @[Mux.scala 27:72]
  wire [1:0] _T_22133 = _T_22792 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22388 = _T_22387 | _T_22133; // @[Mux.scala 27:72]
  wire [1:0] _T_22134 = _T_22794 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22389 = _T_22388 | _T_22134; // @[Mux.scala 27:72]
  wire [1:0] _T_22135 = _T_22796 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22390 = _T_22389 | _T_22135; // @[Mux.scala 27:72]
  wire [1:0] _T_22136 = _T_22798 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22391 = _T_22390 | _T_22136; // @[Mux.scala 27:72]
  wire [1:0] _T_22137 = _T_22800 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22392 = _T_22391 | _T_22137; // @[Mux.scala 27:72]
  wire [1:0] _T_22138 = _T_22802 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22393 = _T_22392 | _T_22138; // @[Mux.scala 27:72]
  wire [1:0] _T_22139 = _T_22804 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22394 = _T_22393 | _T_22139; // @[Mux.scala 27:72]
  wire [1:0] _T_22140 = _T_22806 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22395 = _T_22394 | _T_22140; // @[Mux.scala 27:72]
  wire [1:0] _T_22141 = _T_22808 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22396 = _T_22395 | _T_22141; // @[Mux.scala 27:72]
  wire [1:0] _T_22142 = _T_22810 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22397 = _T_22396 | _T_22142; // @[Mux.scala 27:72]
  wire [1:0] _T_22143 = _T_22812 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22398 = _T_22397 | _T_22143; // @[Mux.scala 27:72]
  wire [1:0] _T_22144 = _T_22814 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22399 = _T_22398 | _T_22144; // @[Mux.scala 27:72]
  wire [1:0] _T_22145 = _T_22816 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22400 = _T_22399 | _T_22145; // @[Mux.scala 27:72]
  wire [1:0] _T_22146 = _T_22818 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22401 = _T_22400 | _T_22146; // @[Mux.scala 27:72]
  wire [1:0] _T_22147 = _T_22820 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22402 = _T_22401 | _T_22147; // @[Mux.scala 27:72]
  wire [1:0] _T_22148 = _T_22822 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22403 = _T_22402 | _T_22148; // @[Mux.scala 27:72]
  wire [1:0] _T_22149 = _T_22824 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22404 = _T_22403 | _T_22149; // @[Mux.scala 27:72]
  wire [1:0] _T_22150 = _T_22826 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22405 = _T_22404 | _T_22150; // @[Mux.scala 27:72]
  wire [1:0] _T_22151 = _T_22828 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22406 = _T_22405 | _T_22151; // @[Mux.scala 27:72]
  wire [1:0] _T_22152 = _T_22830 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22407 = _T_22406 | _T_22152; // @[Mux.scala 27:72]
  wire [1:0] _T_22153 = _T_22832 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22408 = _T_22407 | _T_22153; // @[Mux.scala 27:72]
  wire [1:0] _T_22154 = _T_22834 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22409 = _T_22408 | _T_22154; // @[Mux.scala 27:72]
  wire [1:0] _T_22155 = _T_22836 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22410 = _T_22409 | _T_22155; // @[Mux.scala 27:72]
  wire [1:0] _T_22156 = _T_22838 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22411 = _T_22410 | _T_22156; // @[Mux.scala 27:72]
  wire [1:0] _T_22157 = _T_22840 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22412 = _T_22411 | _T_22157; // @[Mux.scala 27:72]
  wire [1:0] _T_22158 = _T_22842 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22413 = _T_22412 | _T_22158; // @[Mux.scala 27:72]
  wire [1:0] _T_22159 = _T_22844 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22414 = _T_22413 | _T_22159; // @[Mux.scala 27:72]
  wire [1:0] _T_22160 = _T_22846 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22415 = _T_22414 | _T_22160; // @[Mux.scala 27:72]
  wire [1:0] _T_22161 = _T_22848 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22416 = _T_22415 | _T_22161; // @[Mux.scala 27:72]
  wire [1:0] _T_22162 = _T_22850 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22417 = _T_22416 | _T_22162; // @[Mux.scala 27:72]
  wire [1:0] _T_22163 = _T_22852 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22418 = _T_22417 | _T_22163; // @[Mux.scala 27:72]
  wire [1:0] _T_22164 = _T_22854 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22419 = _T_22418 | _T_22164; // @[Mux.scala 27:72]
  wire [1:0] _T_22165 = _T_22856 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22420 = _T_22419 | _T_22165; // @[Mux.scala 27:72]
  wire [1:0] _T_22166 = _T_22858 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22421 = _T_22420 | _T_22166; // @[Mux.scala 27:72]
  wire [1:0] _T_22167 = _T_22860 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22422 = _T_22421 | _T_22167; // @[Mux.scala 27:72]
  wire [1:0] _T_22168 = _T_22862 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22423 = _T_22422 | _T_22168; // @[Mux.scala 27:72]
  wire [1:0] _T_22169 = _T_22864 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22424 = _T_22423 | _T_22169; // @[Mux.scala 27:72]
  wire [1:0] _T_22170 = _T_22866 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22425 = _T_22424 | _T_22170; // @[Mux.scala 27:72]
  wire [1:0] _T_22171 = _T_22868 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22426 = _T_22425 | _T_22171; // @[Mux.scala 27:72]
  wire [1:0] _T_22172 = _T_22870 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22427 = _T_22426 | _T_22172; // @[Mux.scala 27:72]
  wire [1:0] _T_22173 = _T_22872 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22428 = _T_22427 | _T_22173; // @[Mux.scala 27:72]
  wire [1:0] _T_22174 = _T_22874 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22429 = _T_22428 | _T_22174; // @[Mux.scala 27:72]
  wire [1:0] _T_22175 = _T_22876 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22430 = _T_22429 | _T_22175; // @[Mux.scala 27:72]
  wire [1:0] _T_22176 = _T_22878 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22431 = _T_22430 | _T_22176; // @[Mux.scala 27:72]
  wire [1:0] _T_22177 = _T_22880 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22432 = _T_22431 | _T_22177; // @[Mux.scala 27:72]
  wire [1:0] _T_22178 = _T_22882 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22433 = _T_22432 | _T_22178; // @[Mux.scala 27:72]
  wire [1:0] _T_22179 = _T_22884 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22434 = _T_22433 | _T_22179; // @[Mux.scala 27:72]
  wire [1:0] _T_22180 = _T_22886 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22435 = _T_22434 | _T_22180; // @[Mux.scala 27:72]
  wire [1:0] _T_22181 = _T_22888 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22436 = _T_22435 | _T_22181; // @[Mux.scala 27:72]
  wire [1:0] _T_22182 = _T_22890 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22437 = _T_22436 | _T_22182; // @[Mux.scala 27:72]
  wire [1:0] _T_22183 = _T_22892 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22438 = _T_22437 | _T_22183; // @[Mux.scala 27:72]
  wire [1:0] _T_22184 = _T_22894 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22439 = _T_22438 | _T_22184; // @[Mux.scala 27:72]
  wire [1:0] _T_22185 = _T_22896 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22440 = _T_22439 | _T_22185; // @[Mux.scala 27:72]
  wire [1:0] _T_22186 = _T_22898 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22441 = _T_22440 | _T_22186; // @[Mux.scala 27:72]
  wire [1:0] _T_22187 = _T_22900 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22442 = _T_22441 | _T_22187; // @[Mux.scala 27:72]
  wire [1:0] _T_22188 = _T_22902 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22443 = _T_22442 | _T_22188; // @[Mux.scala 27:72]
  wire [1:0] _T_22189 = _T_22904 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22444 = _T_22443 | _T_22189; // @[Mux.scala 27:72]
  wire [1:0] _T_22190 = _T_22906 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22445 = _T_22444 | _T_22190; // @[Mux.scala 27:72]
  wire [1:0] _T_22191 = _T_22908 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22446 = _T_22445 | _T_22191; // @[Mux.scala 27:72]
  wire [1:0] _T_22192 = _T_22910 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22447 = _T_22446 | _T_22192; // @[Mux.scala 27:72]
  wire [1:0] _T_22193 = _T_22912 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22448 = _T_22447 | _T_22193; // @[Mux.scala 27:72]
  wire [1:0] _T_22194 = _T_22914 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22449 = _T_22448 | _T_22194; // @[Mux.scala 27:72]
  wire [1:0] _T_22195 = _T_22916 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22450 = _T_22449 | _T_22195; // @[Mux.scala 27:72]
  wire [1:0] _T_22196 = _T_22918 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22451 = _T_22450 | _T_22196; // @[Mux.scala 27:72]
  wire [1:0] _T_22197 = _T_22920 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22452 = _T_22451 | _T_22197; // @[Mux.scala 27:72]
  wire [1:0] _T_22198 = _T_22922 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22453 = _T_22452 | _T_22198; // @[Mux.scala 27:72]
  wire [1:0] _T_22199 = _T_22924 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22454 = _T_22453 | _T_22199; // @[Mux.scala 27:72]
  wire [1:0] _T_22200 = _T_22926 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22455 = _T_22454 | _T_22200; // @[Mux.scala 27:72]
  wire [1:0] _T_22201 = _T_22928 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22456 = _T_22455 | _T_22201; // @[Mux.scala 27:72]
  wire [1:0] _T_22202 = _T_22930 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22457 = _T_22456 | _T_22202; // @[Mux.scala 27:72]
  wire [1:0] _T_22203 = _T_22932 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22458 = _T_22457 | _T_22203; // @[Mux.scala 27:72]
  wire [1:0] _T_22204 = _T_22934 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22459 = _T_22458 | _T_22204; // @[Mux.scala 27:72]
  wire [1:0] _T_22205 = _T_22936 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22460 = _T_22459 | _T_22205; // @[Mux.scala 27:72]
  wire [1:0] _T_22206 = _T_22938 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22461 = _T_22460 | _T_22206; // @[Mux.scala 27:72]
  wire [1:0] _T_22207 = _T_22940 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22462 = _T_22461 | _T_22207; // @[Mux.scala 27:72]
  wire [1:0] _T_22208 = _T_22942 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22463 = _T_22462 | _T_22208; // @[Mux.scala 27:72]
  wire [1:0] _T_22209 = _T_22944 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22464 = _T_22463 | _T_22209; // @[Mux.scala 27:72]
  wire [1:0] _T_22210 = _T_22946 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22465 = _T_22464 | _T_22210; // @[Mux.scala 27:72]
  wire [1:0] _T_22211 = _T_22948 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22466 = _T_22465 | _T_22211; // @[Mux.scala 27:72]
  wire [1:0] _T_22212 = _T_22950 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22467 = _T_22466 | _T_22212; // @[Mux.scala 27:72]
  wire [1:0] _T_22213 = _T_22952 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22468 = _T_22467 | _T_22213; // @[Mux.scala 27:72]
  wire [1:0] _T_22214 = _T_22954 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22469 = _T_22468 | _T_22214; // @[Mux.scala 27:72]
  wire [1:0] _T_22215 = _T_22956 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22470 = _T_22469 | _T_22215; // @[Mux.scala 27:72]
  wire [1:0] _T_22216 = _T_22958 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22471 = _T_22470 | _T_22216; // @[Mux.scala 27:72]
  wire [1:0] _T_22217 = _T_22960 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22472 = _T_22471 | _T_22217; // @[Mux.scala 27:72]
  wire [1:0] _T_22218 = _T_22962 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22473 = _T_22472 | _T_22218; // @[Mux.scala 27:72]
  wire [1:0] _T_22219 = _T_22964 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22474 = _T_22473 | _T_22219; // @[Mux.scala 27:72]
  wire [1:0] _T_22220 = _T_22966 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22475 = _T_22474 | _T_22220; // @[Mux.scala 27:72]
  wire [1:0] _T_22221 = _T_22968 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22476 = _T_22475 | _T_22221; // @[Mux.scala 27:72]
  wire [1:0] _T_22222 = _T_22970 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22477 = _T_22476 | _T_22222; // @[Mux.scala 27:72]
  wire [1:0] _T_22223 = _T_22972 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22478 = _T_22477 | _T_22223; // @[Mux.scala 27:72]
  wire [1:0] _T_22224 = _T_22974 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22479 = _T_22478 | _T_22224; // @[Mux.scala 27:72]
  wire [1:0] _T_22225 = _T_22976 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22480 = _T_22479 | _T_22225; // @[Mux.scala 27:72]
  wire [1:0] _T_22226 = _T_22978 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22481 = _T_22480 | _T_22226; // @[Mux.scala 27:72]
  wire [1:0] _T_22227 = _T_22980 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22482 = _T_22481 | _T_22227; // @[Mux.scala 27:72]
  wire [1:0] _T_22228 = _T_22982 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22483 = _T_22482 | _T_22228; // @[Mux.scala 27:72]
  wire [1:0] _T_22229 = _T_22984 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22484 = _T_22483 | _T_22229; // @[Mux.scala 27:72]
  wire [1:0] _T_22230 = _T_22986 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22485 = _T_22484 | _T_22230; // @[Mux.scala 27:72]
  wire [1:0] _T_22231 = _T_22988 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22486 = _T_22485 | _T_22231; // @[Mux.scala 27:72]
  wire [1:0] _T_22232 = _T_22990 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22487 = _T_22486 | _T_22232; // @[Mux.scala 27:72]
  wire [1:0] _T_22233 = _T_22992 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22488 = _T_22487 | _T_22233; // @[Mux.scala 27:72]
  wire [1:0] _T_22234 = _T_22994 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22489 = _T_22488 | _T_22234; // @[Mux.scala 27:72]
  wire [1:0] _T_22235 = _T_22996 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22490 = _T_22489 | _T_22235; // @[Mux.scala 27:72]
  wire [1:0] _T_22236 = _T_22998 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22491 = _T_22490 | _T_22236; // @[Mux.scala 27:72]
  wire [1:0] _T_22237 = _T_23000 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22492 = _T_22491 | _T_22237; // @[Mux.scala 27:72]
  wire [1:0] _T_22238 = _T_23002 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22493 = _T_22492 | _T_22238; // @[Mux.scala 27:72]
  wire [1:0] _T_22239 = _T_23004 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22494 = _T_22493 | _T_22239; // @[Mux.scala 27:72]
  wire [1:0] _T_22240 = _T_23006 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22495 = _T_22494 | _T_22240; // @[Mux.scala 27:72]
  wire [1:0] _T_22241 = _T_23008 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_f = _T_22495 | _T_22241; // @[Mux.scala 27:72]
  wire [1:0] _T_271 = _T_162 ? bht_bank0_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_272 = io_ifc_fetch_addr_f[0] ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank0_rd_data_f = _T_271 | _T_272; // @[Mux.scala 27:72]
  wire  _T_289 = bht_force_taken_f[0] | bht_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 299:45]
  wire  _T_291 = _T_289 & bht_valid_f[0]; // @[ifu_bp_ctl.scala 299:72]
  wire [1:0] bht_dir_f = {_T_286,_T_291}; // @[Cat.scala 29:58]
  wire  _T_14 = ~bht_dir_f[0]; // @[ifu_bp_ctl.scala 119:23]
  wire [1:0] btb_sel_f = {_T_14,bht_dir_f[0]}; // @[Cat.scala 29:58]
  wire [1:0] fetch_start_f = {io_ifc_fetch_addr_f[0],_T_162}; // @[Cat.scala 29:58]
  wire  _T_38 = io_exu_bp_exu_mp_btag == _T_30; // @[ifu_bp_ctl.scala 140:53]
  wire  _T_39 = _T_38 & exu_mp_valid; // @[ifu_bp_ctl.scala 140:73]
  wire  _T_40 = _T_39 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 140:88]
  wire  _T_41 = io_exu_bp_exu_mp_index == btb_rd_addr_f; // @[ifu_bp_ctl.scala 140:124]
  wire  _T_42 = _T_40 & _T_41; // @[ifu_bp_ctl.scala 140:109]
  wire  _T_43 = io_exu_bp_exu_mp_btag == _T_37; // @[ifu_bp_ctl.scala 141:56]
  wire  _T_44 = _T_43 & exu_mp_valid; // @[ifu_bp_ctl.scala 141:79]
  wire  _T_45 = _T_44 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 141:94]
  wire  _T_46 = io_exu_bp_exu_mp_index == btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 141:130]
  wire  _T_47 = _T_45 & _T_46; // @[ifu_bp_ctl.scala 141:115]
  wire [1:0] _T_168 = ~bht_valid_f; // @[ifu_bp_ctl.scala 194:44]
  reg  exu_mp_way_f; // @[Reg.scala 27:20]
  wire [255:0] _T_172 = 256'h1 << btb_rd_addr_f; // @[ifu_bp_ctl.scala 213:31]
  reg [255:0] btb_lru_b0_f; // @[Reg.scala 27:20]
  wire [255:0] _T_205 = _T_172 & btb_lru_b0_f; // @[ifu_bp_ctl.scala 239:78]
  wire  _T_206 = |_T_205; // @[ifu_bp_ctl.scala 239:94]
  wire  _T_207 = _T_42 ? exu_mp_way_f : _T_206; // @[ifu_bp_ctl.scala 239:25]
  wire [1:0] _T_214 = {_T_207,_T_207}; // @[Cat.scala 29:58]
  wire [1:0] _T_218 = _T_162 ? _T_214 : 2'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_173 = 256'h1 << btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 216:34]
  wire [255:0] _T_209 = _T_173 & btb_lru_b0_f; // @[ifu_bp_ctl.scala 241:87]
  wire  _T_210 = |_T_209; // @[ifu_bp_ctl.scala 241:103]
  wire  _T_211 = _T_47 ? exu_mp_way_f : _T_210; // @[ifu_bp_ctl.scala 241:28]
  wire [1:0] _T_217 = {_T_211,_T_207}; // @[Cat.scala 29:58]
  wire [1:0] _T_219 = io_ifc_fetch_addr_f[0] ? _T_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] btb_vlru_rd_f = _T_218 | _T_219; // @[Mux.scala 27:72]
  wire [1:0] _T_169 = _T_168 & btb_vlru_rd_f; // @[ifu_bp_ctl.scala 194:55]
  wire [1:0] _T_230 = _T_162 ? _T_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_229 = {_T_127[0],_T_107[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_231 = io_ifc_fetch_addr_f[0] ? _T_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] tag_match_vway1_expanded_f = _T_230 | _T_231; // @[Mux.scala 27:72]
  wire [255:0] _T_171 = 256'h1 << io_exu_bp_exu_mp_index; // @[ifu_bp_ctl.scala 210:28]
  wire [255:0] _T_175 = exu_mp_valid ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] _T_176 = _T_171 & _T_175; // @[ifu_bp_ctl.scala 219:36]
  wire  _T_179 = bht_valid_f[0] | bht_valid_f[1]; // @[ifu_bp_ctl.scala 222:42]
  wire  _T_180 = _T_179 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 222:58]
  wire  _T_182 = _T_180 & _T; // @[ifu_bp_ctl.scala 222:79]
  wire [255:0] _T_184 = _T_182 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] _T_185 = _T_172 & _T_184; // @[ifu_bp_ctl.scala 224:42]
  wire [255:0] _T_188 = _T_173 & _T_184; // @[ifu_bp_ctl.scala 225:48]
  wire [255:0] _T_189 = ~_T_176; // @[ifu_bp_ctl.scala 227:25]
  wire [255:0] _T_190 = ~_T_185; // @[ifu_bp_ctl.scala 227:40]
  wire [255:0] _T_191 = _T_189 & _T_190; // @[ifu_bp_ctl.scala 227:38]
  wire  _T_193 = ~io_exu_bp_exu_mp_pkt_bits_way; // @[ifu_bp_ctl.scala 234:39]
  wire [255:0] _T_196 = _T_193 ? _T_176 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_197 = _T_57 ? _T_185 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_198 = _T_77 ? _T_188 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_199 = _T_196 | _T_197; // @[Mux.scala 27:72]
  wire [255:0] _T_200 = _T_199 | _T_198; // @[Mux.scala 27:72]
  wire [255:0] _T_202 = _T_191 & btb_lru_b0_f; // @[ifu_bp_ctl.scala 236:73]
  wire [255:0] _T_203 = _T_200 | _T_202; // @[ifu_bp_ctl.scala 236:55]
  wire  _T_234 = io_ifc_fetch_req_f | exu_mp_valid; // @[ifu_bp_ctl.scala 251:60]
  wire [15:0] _T_249 = btb_sel_f[1] ? btb_vbank1_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_250 = btb_sel_f[0] ? btb_vbank0_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] btb_sel_data_f = _T_249 | _T_250; // @[Mux.scala 27:72]
  wire [11:0] btb_rd_tgt_f = btb_sel_data_f[15:4]; // @[ifu_bp_ctl.scala 267:36]
  wire  btb_rd_pc4_f = btb_sel_data_f[3]; // @[ifu_bp_ctl.scala 268:36]
  wire  btb_rd_call_f = btb_sel_data_f[1]; // @[ifu_bp_ctl.scala 269:37]
  wire  btb_rd_ret_f = btb_sel_data_f[0]; // @[ifu_bp_ctl.scala 270:36]
  wire [1:0] _T_299 = {bht_vbank1_rd_data_f[1],bht_vbank0_rd_data_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] hist1_raw = bht_force_taken_f | _T_299; // @[ifu_bp_ctl.scala 305:34]
  wire [1:0] _T_253 = bht_valid_f & hist1_raw; // @[ifu_bp_ctl.scala 277:39]
  wire  _T_254 = |_T_253; // @[ifu_bp_ctl.scala 277:52]
  wire  _T_255 = _T_254 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 277:56]
  wire  _T_256 = ~leak_one_f_d1; // @[ifu_bp_ctl.scala 277:79]
  wire  _T_257 = _T_255 & _T_256; // @[ifu_bp_ctl.scala 277:77]
  wire  _T_258 = ~io_dec_bp_dec_tlu_bpred_disable; // @[ifu_bp_ctl.scala 277:96]
  wire  _T_294 = io_ifu_bp_hit_taken_f & btb_sel_f[1]; // @[ifu_bp_ctl.scala 302:51]
  wire  _T_295 = ~io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 302:69]
  wire  _T_305 = bht_valid_f[1] & btb_vbank1_rd_data_f[4]; // @[ifu_bp_ctl.scala 311:34]
  wire  _T_308 = bht_valid_f[0] & btb_vbank0_rd_data_f[4]; // @[ifu_bp_ctl.scala 312:34]
  wire  _T_311 = ~btb_vbank1_rd_data_f[2]; // @[ifu_bp_ctl.scala 315:37]
  wire  _T_312 = bht_valid_f[1] & _T_311; // @[ifu_bp_ctl.scala 315:35]
  wire  _T_314 = _T_312 & btb_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 315:65]
  wire  _T_317 = ~btb_vbank0_rd_data_f[2]; // @[ifu_bp_ctl.scala 316:37]
  wire  _T_318 = bht_valid_f[0] & _T_317; // @[ifu_bp_ctl.scala 316:35]
  wire  _T_320 = _T_318 & btb_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 316:65]
  wire [1:0] num_valids = bht_valid_f[1] + bht_valid_f[0]; // @[ifu_bp_ctl.scala 319:35]
  wire [1:0] _T_323 = btb_sel_f & bht_dir_f; // @[ifu_bp_ctl.scala 322:28]
  wire  final_h = |_T_323; // @[ifu_bp_ctl.scala 322:41]
  wire  _T_324 = num_valids == 2'h2; // @[ifu_bp_ctl.scala 326:41]
  wire [7:0] _T_328 = {fghr[5:0],1'h0,final_h}; // @[Cat.scala 29:58]
  wire  _T_329 = num_valids == 2'h1; // @[ifu_bp_ctl.scala 327:41]
  wire [7:0] _T_332 = {fghr[6:0],final_h}; // @[Cat.scala 29:58]
  wire  _T_333 = num_valids == 2'h0; // @[ifu_bp_ctl.scala 328:41]
  wire [7:0] _T_336 = _T_324 ? _T_328 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_337 = _T_329 ? _T_332 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_338 = _T_333 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_339 = _T_336 | _T_337; // @[Mux.scala 27:72]
  wire [7:0] merged_ghr = _T_339 | _T_338; // @[Mux.scala 27:72]
  reg  exu_flush_final_d1; // @[Reg.scala 27:20]
  wire  _T_342 = ~exu_flush_final_d1; // @[ifu_bp_ctl.scala 337:27]
  wire  _T_343 = _T_342 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 337:47]
  wire  _T_344 = _T_343 & io_ic_hit_f; // @[ifu_bp_ctl.scala 337:70]
  wire  _T_346 = _T_344 & _T_256; // @[ifu_bp_ctl.scala 337:84]
  wire  _T_349 = io_ifc_fetch_req_f & io_ic_hit_f; // @[ifu_bp_ctl.scala 338:70]
  wire  _T_351 = _T_349 & _T_256; // @[ifu_bp_ctl.scala 338:84]
  wire  _T_352 = ~_T_351; // @[ifu_bp_ctl.scala 338:49]
  wire  _T_353 = _T_342 & _T_352; // @[ifu_bp_ctl.scala 338:47]
  wire [7:0] _T_355 = exu_flush_final_d1 ? io_exu_bp_exu_mp_fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_356 = _T_346 ? merged_ghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_357 = _T_353 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_358 = _T_355 | _T_356; // @[Mux.scala 27:72]
  wire [7:0] fghr_ns = _T_358 | _T_357; // @[Mux.scala 27:72]
  wire  _T_362 = leak_one_f ^ leak_one_f_d1; // @[lib.scala 453:21]
  wire  _T_363 = |_T_362; // @[lib.scala 453:29]
  wire  _T_366 = io_exu_bp_exu_mp_pkt_bits_way ^ exu_mp_way_f; // @[lib.scala 453:21]
  wire  _T_367 = |_T_366; // @[lib.scala 453:29]
  wire  _T_370 = io_exu_flush_final ^ exu_flush_final_d1; // @[lib.scala 475:21]
  wire  _T_371 = |_T_370; // @[lib.scala 475:29]
  wire [7:0] _T_374 = fghr_ns ^ fghr; // @[lib.scala 453:21]
  wire  _T_375 = |_T_374; // @[lib.scala 453:29]
  wire [1:0] _T_378 = io_dec_bp_dec_tlu_bpred_disable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_379 = ~_T_378; // @[ifu_bp_ctl.scala 350:36]
  wire  _T_383 = ~fetch_start_f[0]; // @[ifu_bp_ctl.scala 354:36]
  wire  _T_384 = bht_dir_f[0] & _T_383; // @[ifu_bp_ctl.scala 354:34]
  wire  _T_388 = _T_14 & fetch_start_f[0]; // @[ifu_bp_ctl.scala 354:72]
  wire  _T_389 = _T_384 | _T_388; // @[ifu_bp_ctl.scala 354:55]
  wire  _T_392 = bht_dir_f[0] & fetch_start_f[0]; // @[ifu_bp_ctl.scala 355:34]
  wire  _T_397 = _T_14 & _T_383; // @[ifu_bp_ctl.scala 355:71]
  wire  _T_398 = _T_392 | _T_397; // @[ifu_bp_ctl.scala 355:54]
  wire [1:0] bloc_f = {_T_389,_T_398}; // @[Cat.scala 29:58]
  wire  _T_402 = _T_14 & io_ifc_fetch_addr_f[0]; // @[ifu_bp_ctl.scala 357:35]
  wire  _T_403 = ~btb_rd_pc4_f; // @[ifu_bp_ctl.scala 357:62]
  wire  use_fa_plus = _T_402 & _T_403; // @[ifu_bp_ctl.scala 357:60]
  wire  _T_406 = fetch_start_f[0] & btb_sel_f[0]; // @[ifu_bp_ctl.scala 359:44]
  wire  btb_fg_crossing_f = _T_406 & btb_rd_pc4_f; // @[ifu_bp_ctl.scala 359:59]
  wire  bp_total_branch_offset_f = bloc_f[1] ^ btb_rd_pc4_f; // @[ifu_bp_ctl.scala 360:43]
  wire  _T_410 = io_ifc_fetch_req_f & _T_295; // @[ifu_bp_ctl.scala 361:117]
  wire  _T_411 = _T_410 & io_ic_hit_f; // @[ifu_bp_ctl.scala 361:142]
  reg [29:0] ifc_fetch_adder_prior; // @[Reg.scala 27:20]
  wire  _T_416 = ~btb_fg_crossing_f; // @[ifu_bp_ctl.scala 366:32]
  wire  _T_417 = ~use_fa_plus; // @[ifu_bp_ctl.scala 366:53]
  wire  _T_418 = _T_416 & _T_417; // @[ifu_bp_ctl.scala 366:51]
  wire [29:0] _T_421 = use_fa_plus ? fetch_addr_p1_f : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_422 = btb_fg_crossing_f ? ifc_fetch_adder_prior : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_423 = _T_418 ? io_ifc_fetch_addr_f[30:1] : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_424 = _T_421 | _T_422; // @[Mux.scala 27:72]
  wire [29:0] adder_pc_in_f = _T_424 | _T_423; // @[Mux.scala 27:72]
  wire [31:0] _T_428 = {adder_pc_in_f,bp_total_branch_offset_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_429 = {btb_rd_tgt_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_432 = _T_428[12:1] + _T_429[12:1]; // @[lib.scala 68:31]
  wire [18:0] _T_435 = _T_428[31:13] + 19'h1; // @[lib.scala 69:27]
  wire [18:0] _T_438 = _T_428[31:13] - 19'h1; // @[lib.scala 70:27]
  wire  _T_441 = ~_T_432[12]; // @[lib.scala 72:28]
  wire  _T_442 = _T_429[12] ^ _T_441; // @[lib.scala 72:26]
  wire  _T_445 = ~_T_429[12]; // @[lib.scala 73:20]
  wire  _T_447 = _T_445 & _T_432[12]; // @[lib.scala 73:26]
  wire  _T_451 = _T_429[12] & _T_441; // @[lib.scala 74:26]
  wire [18:0] _T_453 = _T_442 ? _T_428[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_454 = _T_447 ? _T_435 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_455 = _T_451 ? _T_438 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_456 = _T_453 | _T_454; // @[Mux.scala 27:72]
  wire [18:0] _T_457 = _T_456 | _T_455; // @[Mux.scala 27:72]
  wire [31:0] bp_btb_target_adder_f = {_T_457,_T_432[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_461 = ~btb_rd_call_f; // @[ifu_bp_ctl.scala 374:55]
  wire  _T_462 = btb_rd_ret_f & _T_461; // @[ifu_bp_ctl.scala 374:53]
  reg [31:0] rets_out_0; // @[Reg.scala 27:20]
  wire  _T_464 = _T_462 & rets_out_0[0]; // @[ifu_bp_ctl.scala 374:70]
  wire  _T_465 = _T_464 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 374:87]
  wire [30:0] _T_467 = _T_465 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [30:0] _T_469 = _T_467 & rets_out_0[31:1]; // @[ifu_bp_ctl.scala 374:113]
  wire  _T_474 = ~_T_464; // @[ifu_bp_ctl.scala 375:15]
  wire  _T_475 = _T_474 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 375:65]
  wire [30:0] _T_477 = _T_475 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [30:0] _T_479 = _T_477 & bp_btb_target_adder_f[31:1]; // @[ifu_bp_ctl.scala 375:91]
  wire [12:0] _T_487 = {11'h0,_T_403,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_490 = _T_428[12:1] + _T_487[12:1]; // @[lib.scala 68:31]
  wire  _T_499 = ~_T_490[12]; // @[lib.scala 72:28]
  wire  _T_500 = _T_487[12] ^ _T_499; // @[lib.scala 72:26]
  wire  _T_503 = ~_T_487[12]; // @[lib.scala 73:20]
  wire  _T_505 = _T_503 & _T_490[12]; // @[lib.scala 73:26]
  wire  _T_509 = _T_487[12] & _T_499; // @[lib.scala 74:26]
  wire [18:0] _T_511 = _T_500 ? _T_428[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_512 = _T_505 ? _T_435 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_513 = _T_509 ? _T_438 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_514 = _T_511 | _T_512; // @[Mux.scala 27:72]
  wire [18:0] _T_515 = _T_514 | _T_513; // @[Mux.scala 27:72]
  wire [31:0] bp_rs_call_target_f = {_T_515,_T_490[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_519 = ~btb_rd_ret_f; // @[ifu_bp_ctl.scala 379:33]
  wire  _T_520 = btb_rd_call_f & _T_519; // @[ifu_bp_ctl.scala 379:31]
  wire  rs_push = _T_520 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 379:47]
  wire  rs_pop = _T_462 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 380:46]
  wire  _T_523 = ~rs_push; // @[ifu_bp_ctl.scala 381:17]
  wire  _T_524 = ~rs_pop; // @[ifu_bp_ctl.scala 381:28]
  wire  rs_hold = _T_523 & _T_524; // @[ifu_bp_ctl.scala 381:26]
  wire  rsenable_0 = ~rs_hold; // @[ifu_bp_ctl.scala 383:60]
  wire  rsenable_1 = rs_push | rs_pop; // @[ifu_bp_ctl.scala 383:119]
  wire [31:0] _T_527 = {bp_rs_call_target_f[31:1],1'h1}; // @[Cat.scala 29:58]
  wire [31:0] _T_529 = rs_push ? _T_527 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_1; // @[Reg.scala 27:20]
  wire [31:0] _T_530 = rs_pop ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_0 = _T_529 | _T_530; // @[Mux.scala 27:72]
  wire [31:0] _T_534 = rs_push ? rets_out_0 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_2; // @[Reg.scala 27:20]
  wire [31:0] _T_535 = rs_pop ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_1 = _T_534 | _T_535; // @[Mux.scala 27:72]
  wire [31:0] _T_539 = rs_push ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_3; // @[Reg.scala 27:20]
  wire [31:0] _T_540 = rs_pop ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_2 = _T_539 | _T_540; // @[Mux.scala 27:72]
  wire [31:0] _T_544 = rs_push ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_4; // @[Reg.scala 27:20]
  wire [31:0] _T_545 = rs_pop ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_3 = _T_544 | _T_545; // @[Mux.scala 27:72]
  wire [31:0] _T_549 = rs_push ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_5; // @[Reg.scala 27:20]
  wire [31:0] _T_550 = rs_pop ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_4 = _T_549 | _T_550; // @[Mux.scala 27:72]
  wire [31:0] _T_554 = rs_push ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_6; // @[Reg.scala 27:20]
  wire [31:0] _T_555 = rs_pop ? rets_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_5 = _T_554 | _T_555; // @[Mux.scala 27:72]
  wire [31:0] _T_559 = rs_push ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_7; // @[Reg.scala 27:20]
  wire [31:0] _T_560 = rs_pop ? rets_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_6 = _T_559 | _T_560; // @[Mux.scala 27:72]
  wire  _T_578 = ~dec_tlu_error_wb; // @[ifu_bp_ctl.scala 395:35]
  wire  btb_valid = exu_mp_valid & _T_578; // @[ifu_bp_ctl.scala 395:32]
  wire  _T_579 = io_exu_bp_exu_mp_pkt_bits_pcall | io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 399:89]
  wire  _T_580 = io_exu_bp_exu_mp_pkt_bits_pret | io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 399:113]
  wire [21:0] btb_wr_data = {io_exu_bp_exu_mp_btag,io_exu_bp_exu_mp_pkt_bits_toffset,io_exu_bp_exu_mp_pkt_bits_pc4,io_exu_bp_exu_mp_pkt_bits_boffset,_T_579,_T_580,btb_valid}; // @[Cat.scala 29:58]
  wire  _T_586 = exu_mp_valid & io_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu_bp_ctl.scala 400:41]
  wire  _T_587 = ~io_exu_bp_exu_mp_pkt_valid; // @[ifu_bp_ctl.scala 400:59]
  wire  exu_mp_valid_write = _T_586 & _T_587; // @[ifu_bp_ctl.scala 400:57]
  wire  middle_of_bank = io_exu_bp_exu_mp_pkt_bits_pc4 ^ io_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu_bp_ctl.scala 401:35]
  wire  _T_588 = ~io_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu_bp_ctl.scala 404:43]
  wire  _T_589 = exu_mp_valid & _T_588; // @[ifu_bp_ctl.scala 404:41]
  wire  _T_590 = ~io_exu_bp_exu_mp_pkt_bits_pret; // @[ifu_bp_ctl.scala 404:58]
  wire  _T_591 = _T_589 & _T_590; // @[ifu_bp_ctl.scala 404:56]
  wire  _T_592 = ~io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 404:72]
  wire  _T_593 = _T_591 & _T_592; // @[ifu_bp_ctl.scala 404:70]
  wire [1:0] _T_595 = _T_593 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_596 = ~middle_of_bank; // @[ifu_bp_ctl.scala 404:106]
  wire [1:0] _T_597 = {middle_of_bank,_T_596}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en0 = _T_595 & _T_597; // @[ifu_bp_ctl.scala 404:84]
  wire [1:0] _T_599 = io_dec_bp_dec_tlu_br0_r_pkt_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_600 = ~io_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu_bp_ctl.scala 405:75]
  wire [1:0] _T_601 = {io_dec_bp_dec_tlu_br0_r_pkt_bits_middle,_T_600}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en2 = _T_599 & _T_601; // @[ifu_bp_ctl.scala 405:46]
  wire [9:0] _T_602 = {io_exu_bp_exu_mp_index,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_wr_addr0 = _T_602[9:2] ^ io_exu_bp_exu_mp_eghr; // @[lib.scala 56:35]
  wire [9:0] _T_605 = {io_exu_bp_exu_i0_br_index_r,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_wr_addr2 = _T_605[9:2] ^ io_exu_bp_exu_i0_br_fghr_r; // @[lib.scala 56:35]
  wire  _T_615 = _T_193 & exu_mp_valid_write; // @[ifu_bp_ctl.scala 424:39]
  wire  _T_617 = _T_615 & _T_578; // @[ifu_bp_ctl.scala 424:60]
  wire  _T_618 = ~io_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu_bp_ctl.scala 424:87]
  wire  _T_619 = _T_618 & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 424:104]
  wire  _T_620 = _T_617 | _T_619; // @[ifu_bp_ctl.scala 424:83]
  wire  _T_621 = io_exu_bp_exu_mp_pkt_bits_way & exu_mp_valid_write; // @[ifu_bp_ctl.scala 425:36]
  wire  _T_623 = _T_621 & _T_578; // @[ifu_bp_ctl.scala 425:57]
  wire  _T_624 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 425:98]
  wire  _T_625 = _T_623 | _T_624; // @[ifu_bp_ctl.scala 425:80]
  wire [7:0] _T_627 = dec_tlu_error_wb ? io_exu_bp_exu_i0_br_index_r : io_exu_bp_exu_mp_index; // @[ifu_bp_ctl.scala 428:24]
  wire  _T_642 = _T_627 == 8'h0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_643 = _T_642 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_646 = _T_627 == 8'h1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_647 = _T_646 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_650 = _T_627 == 8'h2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_651 = _T_650 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_654 = _T_627 == 8'h3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_655 = _T_654 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_658 = _T_627 == 8'h4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_659 = _T_658 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_662 = _T_627 == 8'h5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_663 = _T_662 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_666 = _T_627 == 8'h6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_667 = _T_666 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_670 = _T_627 == 8'h7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_671 = _T_670 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_674 = _T_627 == 8'h8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_675 = _T_674 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_678 = _T_627 == 8'h9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_679 = _T_678 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_682 = _T_627 == 8'ha; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_683 = _T_682 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_686 = _T_627 == 8'hb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_687 = _T_686 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_690 = _T_627 == 8'hc; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_691 = _T_690 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_694 = _T_627 == 8'hd; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_695 = _T_694 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_698 = _T_627 == 8'he; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_699 = _T_698 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_702 = _T_627 == 8'hf; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_703 = _T_702 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_706 = _T_627 == 8'h10; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_707 = _T_706 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_710 = _T_627 == 8'h11; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_711 = _T_710 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_714 = _T_627 == 8'h12; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_715 = _T_714 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_718 = _T_627 == 8'h13; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_719 = _T_718 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_722 = _T_627 == 8'h14; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_723 = _T_722 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_726 = _T_627 == 8'h15; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_727 = _T_726 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_730 = _T_627 == 8'h16; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_731 = _T_730 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_734 = _T_627 == 8'h17; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_735 = _T_734 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_738 = _T_627 == 8'h18; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_739 = _T_738 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_742 = _T_627 == 8'h19; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_743 = _T_742 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_746 = _T_627 == 8'h1a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_747 = _T_746 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_750 = _T_627 == 8'h1b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_751 = _T_750 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_754 = _T_627 == 8'h1c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_755 = _T_754 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_758 = _T_627 == 8'h1d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_759 = _T_758 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_762 = _T_627 == 8'h1e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_763 = _T_762 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_766 = _T_627 == 8'h1f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_767 = _T_766 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_770 = _T_627 == 8'h20; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_771 = _T_770 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_774 = _T_627 == 8'h21; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_775 = _T_774 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_778 = _T_627 == 8'h22; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_779 = _T_778 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_782 = _T_627 == 8'h23; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_783 = _T_782 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_786 = _T_627 == 8'h24; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_787 = _T_786 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_790 = _T_627 == 8'h25; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_791 = _T_790 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_794 = _T_627 == 8'h26; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_795 = _T_794 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_798 = _T_627 == 8'h27; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_799 = _T_798 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_802 = _T_627 == 8'h28; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_803 = _T_802 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_806 = _T_627 == 8'h29; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_807 = _T_806 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_810 = _T_627 == 8'h2a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_811 = _T_810 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_814 = _T_627 == 8'h2b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_815 = _T_814 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_818 = _T_627 == 8'h2c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_819 = _T_818 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_822 = _T_627 == 8'h2d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_823 = _T_822 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_826 = _T_627 == 8'h2e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_827 = _T_826 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_830 = _T_627 == 8'h2f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_831 = _T_830 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_834 = _T_627 == 8'h30; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_835 = _T_834 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_838 = _T_627 == 8'h31; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_839 = _T_838 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_842 = _T_627 == 8'h32; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_843 = _T_842 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_846 = _T_627 == 8'h33; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_847 = _T_846 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_850 = _T_627 == 8'h34; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_851 = _T_850 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_854 = _T_627 == 8'h35; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_855 = _T_854 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_858 = _T_627 == 8'h36; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_859 = _T_858 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_862 = _T_627 == 8'h37; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_863 = _T_862 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_866 = _T_627 == 8'h38; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_867 = _T_866 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_870 = _T_627 == 8'h39; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_871 = _T_870 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_874 = _T_627 == 8'h3a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_875 = _T_874 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_878 = _T_627 == 8'h3b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_879 = _T_878 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_882 = _T_627 == 8'h3c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_883 = _T_882 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_886 = _T_627 == 8'h3d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_887 = _T_886 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_890 = _T_627 == 8'h3e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_891 = _T_890 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_894 = _T_627 == 8'h3f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_895 = _T_894 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_898 = _T_627 == 8'h40; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_899 = _T_898 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_902 = _T_627 == 8'h41; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_903 = _T_902 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_906 = _T_627 == 8'h42; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_907 = _T_906 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_910 = _T_627 == 8'h43; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_911 = _T_910 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_914 = _T_627 == 8'h44; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_915 = _T_914 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_918 = _T_627 == 8'h45; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_919 = _T_918 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_922 = _T_627 == 8'h46; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_923 = _T_922 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_926 = _T_627 == 8'h47; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_927 = _T_926 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_930 = _T_627 == 8'h48; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_931 = _T_930 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_934 = _T_627 == 8'h49; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_935 = _T_934 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_938 = _T_627 == 8'h4a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_939 = _T_938 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_942 = _T_627 == 8'h4b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_943 = _T_942 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_946 = _T_627 == 8'h4c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_947 = _T_946 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_950 = _T_627 == 8'h4d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_951 = _T_950 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_954 = _T_627 == 8'h4e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_955 = _T_954 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_958 = _T_627 == 8'h4f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_959 = _T_958 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_962 = _T_627 == 8'h50; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_963 = _T_962 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_966 = _T_627 == 8'h51; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_967 = _T_966 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_970 = _T_627 == 8'h52; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_971 = _T_970 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_974 = _T_627 == 8'h53; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_975 = _T_974 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_978 = _T_627 == 8'h54; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_979 = _T_978 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_982 = _T_627 == 8'h55; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_983 = _T_982 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_986 = _T_627 == 8'h56; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_987 = _T_986 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_990 = _T_627 == 8'h57; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_991 = _T_990 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_994 = _T_627 == 8'h58; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_995 = _T_994 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_998 = _T_627 == 8'h59; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_999 = _T_998 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1002 = _T_627 == 8'h5a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1003 = _T_1002 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1006 = _T_627 == 8'h5b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1007 = _T_1006 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1010 = _T_627 == 8'h5c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1011 = _T_1010 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1014 = _T_627 == 8'h5d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1015 = _T_1014 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1018 = _T_627 == 8'h5e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1019 = _T_1018 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1022 = _T_627 == 8'h5f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1023 = _T_1022 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1026 = _T_627 == 8'h60; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1027 = _T_1026 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1030 = _T_627 == 8'h61; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1031 = _T_1030 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1034 = _T_627 == 8'h62; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1035 = _T_1034 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1038 = _T_627 == 8'h63; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1039 = _T_1038 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1042 = _T_627 == 8'h64; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1043 = _T_1042 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1046 = _T_627 == 8'h65; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1047 = _T_1046 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1050 = _T_627 == 8'h66; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1051 = _T_1050 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1054 = _T_627 == 8'h67; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1055 = _T_1054 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1058 = _T_627 == 8'h68; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1059 = _T_1058 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1062 = _T_627 == 8'h69; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1063 = _T_1062 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1066 = _T_627 == 8'h6a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1067 = _T_1066 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1070 = _T_627 == 8'h6b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1071 = _T_1070 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1074 = _T_627 == 8'h6c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1075 = _T_1074 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1078 = _T_627 == 8'h6d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1079 = _T_1078 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1082 = _T_627 == 8'h6e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1083 = _T_1082 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1086 = _T_627 == 8'h6f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1087 = _T_1086 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1090 = _T_627 == 8'h70; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1091 = _T_1090 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1094 = _T_627 == 8'h71; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1095 = _T_1094 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1098 = _T_627 == 8'h72; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1099 = _T_1098 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1102 = _T_627 == 8'h73; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1103 = _T_1102 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1106 = _T_627 == 8'h74; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1107 = _T_1106 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1110 = _T_627 == 8'h75; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1111 = _T_1110 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1114 = _T_627 == 8'h76; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1115 = _T_1114 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1118 = _T_627 == 8'h77; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1119 = _T_1118 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1122 = _T_627 == 8'h78; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1123 = _T_1122 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1126 = _T_627 == 8'h79; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1127 = _T_1126 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1130 = _T_627 == 8'h7a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1131 = _T_1130 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1134 = _T_627 == 8'h7b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1135 = _T_1134 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1138 = _T_627 == 8'h7c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1139 = _T_1138 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1142 = _T_627 == 8'h7d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1143 = _T_1142 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1146 = _T_627 == 8'h7e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1147 = _T_1146 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1150 = _T_627 == 8'h7f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1151 = _T_1150 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1154 = _T_627 == 8'h80; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1155 = _T_1154 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1158 = _T_627 == 8'h81; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1159 = _T_1158 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1162 = _T_627 == 8'h82; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1163 = _T_1162 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1166 = _T_627 == 8'h83; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1167 = _T_1166 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1170 = _T_627 == 8'h84; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1171 = _T_1170 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1174 = _T_627 == 8'h85; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1175 = _T_1174 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1178 = _T_627 == 8'h86; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1179 = _T_1178 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1182 = _T_627 == 8'h87; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1183 = _T_1182 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1186 = _T_627 == 8'h88; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1187 = _T_1186 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1190 = _T_627 == 8'h89; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1191 = _T_1190 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1194 = _T_627 == 8'h8a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1195 = _T_1194 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1198 = _T_627 == 8'h8b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1199 = _T_1198 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1202 = _T_627 == 8'h8c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1203 = _T_1202 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1206 = _T_627 == 8'h8d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1207 = _T_1206 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1210 = _T_627 == 8'h8e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1211 = _T_1210 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1214 = _T_627 == 8'h8f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1215 = _T_1214 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1218 = _T_627 == 8'h90; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1219 = _T_1218 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1222 = _T_627 == 8'h91; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1223 = _T_1222 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1226 = _T_627 == 8'h92; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1227 = _T_1226 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1230 = _T_627 == 8'h93; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1231 = _T_1230 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1234 = _T_627 == 8'h94; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1235 = _T_1234 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1238 = _T_627 == 8'h95; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1239 = _T_1238 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1242 = _T_627 == 8'h96; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1243 = _T_1242 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1246 = _T_627 == 8'h97; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1247 = _T_1246 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1250 = _T_627 == 8'h98; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1251 = _T_1250 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1254 = _T_627 == 8'h99; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1255 = _T_1254 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1258 = _T_627 == 8'h9a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1259 = _T_1258 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1262 = _T_627 == 8'h9b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1263 = _T_1262 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1266 = _T_627 == 8'h9c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1267 = _T_1266 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1270 = _T_627 == 8'h9d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1271 = _T_1270 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1274 = _T_627 == 8'h9e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1275 = _T_1274 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1278 = _T_627 == 8'h9f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1279 = _T_1278 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1282 = _T_627 == 8'ha0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1283 = _T_1282 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1286 = _T_627 == 8'ha1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1287 = _T_1286 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1290 = _T_627 == 8'ha2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1291 = _T_1290 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1294 = _T_627 == 8'ha3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1295 = _T_1294 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1298 = _T_627 == 8'ha4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1299 = _T_1298 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1302 = _T_627 == 8'ha5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1303 = _T_1302 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1306 = _T_627 == 8'ha6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1307 = _T_1306 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1310 = _T_627 == 8'ha7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1311 = _T_1310 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1314 = _T_627 == 8'ha8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1315 = _T_1314 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1318 = _T_627 == 8'ha9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1319 = _T_1318 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1322 = _T_627 == 8'haa; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1323 = _T_1322 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1326 = _T_627 == 8'hab; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1327 = _T_1326 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1330 = _T_627 == 8'hac; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1331 = _T_1330 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1334 = _T_627 == 8'had; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1335 = _T_1334 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1338 = _T_627 == 8'hae; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1339 = _T_1338 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1342 = _T_627 == 8'haf; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1343 = _T_1342 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1346 = _T_627 == 8'hb0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1347 = _T_1346 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1350 = _T_627 == 8'hb1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1351 = _T_1350 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1354 = _T_627 == 8'hb2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1355 = _T_1354 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1358 = _T_627 == 8'hb3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1359 = _T_1358 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1362 = _T_627 == 8'hb4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1363 = _T_1362 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1366 = _T_627 == 8'hb5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1367 = _T_1366 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1370 = _T_627 == 8'hb6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1371 = _T_1370 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1374 = _T_627 == 8'hb7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1375 = _T_1374 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1378 = _T_627 == 8'hb8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1379 = _T_1378 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1382 = _T_627 == 8'hb9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1383 = _T_1382 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1386 = _T_627 == 8'hba; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1387 = _T_1386 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1390 = _T_627 == 8'hbb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1391 = _T_1390 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1394 = _T_627 == 8'hbc; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1395 = _T_1394 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1398 = _T_627 == 8'hbd; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1399 = _T_1398 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1402 = _T_627 == 8'hbe; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1403 = _T_1402 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1406 = _T_627 == 8'hbf; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1407 = _T_1406 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1410 = _T_627 == 8'hc0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1411 = _T_1410 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1414 = _T_627 == 8'hc1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1415 = _T_1414 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1418 = _T_627 == 8'hc2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1419 = _T_1418 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1422 = _T_627 == 8'hc3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1423 = _T_1422 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1426 = _T_627 == 8'hc4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1427 = _T_1426 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1430 = _T_627 == 8'hc5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1431 = _T_1430 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1434 = _T_627 == 8'hc6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1435 = _T_1434 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1438 = _T_627 == 8'hc7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1439 = _T_1438 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1442 = _T_627 == 8'hc8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1443 = _T_1442 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1446 = _T_627 == 8'hc9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1447 = _T_1446 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1450 = _T_627 == 8'hca; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1451 = _T_1450 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1454 = _T_627 == 8'hcb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1455 = _T_1454 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1458 = _T_627 == 8'hcc; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1459 = _T_1458 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1462 = _T_627 == 8'hcd; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1463 = _T_1462 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1466 = _T_627 == 8'hce; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1467 = _T_1466 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1470 = _T_627 == 8'hcf; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1471 = _T_1470 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1474 = _T_627 == 8'hd0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1475 = _T_1474 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1478 = _T_627 == 8'hd1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1479 = _T_1478 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1482 = _T_627 == 8'hd2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1483 = _T_1482 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1486 = _T_627 == 8'hd3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1487 = _T_1486 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1490 = _T_627 == 8'hd4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1491 = _T_1490 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1494 = _T_627 == 8'hd5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1495 = _T_1494 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1498 = _T_627 == 8'hd6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1499 = _T_1498 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1502 = _T_627 == 8'hd7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1503 = _T_1502 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1506 = _T_627 == 8'hd8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1507 = _T_1506 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1510 = _T_627 == 8'hd9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1511 = _T_1510 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1514 = _T_627 == 8'hda; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1515 = _T_1514 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1518 = _T_627 == 8'hdb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1519 = _T_1518 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1522 = _T_627 == 8'hdc; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1523 = _T_1522 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1526 = _T_627 == 8'hdd; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1527 = _T_1526 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1530 = _T_627 == 8'hde; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1531 = _T_1530 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1534 = _T_627 == 8'hdf; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1535 = _T_1534 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1538 = _T_627 == 8'he0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1539 = _T_1538 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1542 = _T_627 == 8'he1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1543 = _T_1542 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1546 = _T_627 == 8'he2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1547 = _T_1546 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1550 = _T_627 == 8'he3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1551 = _T_1550 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1554 = _T_627 == 8'he4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1555 = _T_1554 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1558 = _T_627 == 8'he5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1559 = _T_1558 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1562 = _T_627 == 8'he6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1563 = _T_1562 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1566 = _T_627 == 8'he7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1567 = _T_1566 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1570 = _T_627 == 8'he8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1571 = _T_1570 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1574 = _T_627 == 8'he9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1575 = _T_1574 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1578 = _T_627 == 8'hea; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1579 = _T_1578 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1582 = _T_627 == 8'heb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1583 = _T_1582 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1586 = _T_627 == 8'hec; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1587 = _T_1586 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1590 = _T_627 == 8'hed; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1591 = _T_1590 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1594 = _T_627 == 8'hee; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1595 = _T_1594 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1598 = _T_627 == 8'hef; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1599 = _T_1598 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1602 = _T_627 == 8'hf0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1603 = _T_1602 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1606 = _T_627 == 8'hf1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1607 = _T_1606 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1610 = _T_627 == 8'hf2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1611 = _T_1610 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1614 = _T_627 == 8'hf3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1615 = _T_1614 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1618 = _T_627 == 8'hf4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1619 = _T_1618 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1622 = _T_627 == 8'hf5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1623 = _T_1622 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1626 = _T_627 == 8'hf6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1627 = _T_1626 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1630 = _T_627 == 8'hf7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1631 = _T_1630 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1634 = _T_627 == 8'hf8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1635 = _T_1634 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1638 = _T_627 == 8'hf9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1639 = _T_1638 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1642 = _T_627 == 8'hfa; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1643 = _T_1642 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1646 = _T_627 == 8'hfb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1647 = _T_1646 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1650 = _T_627 == 8'hfc; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1651 = _T_1650 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1654 = _T_627 == 8'hfd; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1655 = _T_1654 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1658 = _T_627 == 8'hfe; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1659 = _T_1658 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1662 = _T_627 == 8'hff; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1663 = _T_1662 & _T_620; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1667 = _T_642 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1671 = _T_646 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1675 = _T_650 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1679 = _T_654 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1683 = _T_658 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1687 = _T_662 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1691 = _T_666 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1695 = _T_670 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1699 = _T_674 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1703 = _T_678 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1707 = _T_682 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1711 = _T_686 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1715 = _T_690 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1719 = _T_694 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1723 = _T_698 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1727 = _T_702 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1731 = _T_706 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1735 = _T_710 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1739 = _T_714 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1743 = _T_718 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1747 = _T_722 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1751 = _T_726 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1755 = _T_730 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1759 = _T_734 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1763 = _T_738 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1767 = _T_742 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1771 = _T_746 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1775 = _T_750 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1779 = _T_754 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1783 = _T_758 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1787 = _T_762 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1791 = _T_766 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1795 = _T_770 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1799 = _T_774 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1803 = _T_778 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1807 = _T_782 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1811 = _T_786 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1815 = _T_790 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1819 = _T_794 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1823 = _T_798 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1827 = _T_802 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1831 = _T_806 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1835 = _T_810 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1839 = _T_814 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1843 = _T_818 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1847 = _T_822 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1851 = _T_826 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1855 = _T_830 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1859 = _T_834 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1863 = _T_838 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1867 = _T_842 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1871 = _T_846 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1875 = _T_850 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1879 = _T_854 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1883 = _T_858 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1887 = _T_862 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1891 = _T_866 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1895 = _T_870 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1899 = _T_874 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1903 = _T_878 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1907 = _T_882 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1911 = _T_886 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1915 = _T_890 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1919 = _T_894 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1923 = _T_898 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1927 = _T_902 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1931 = _T_906 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1935 = _T_910 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1939 = _T_914 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1943 = _T_918 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1947 = _T_922 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1951 = _T_926 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1955 = _T_930 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1959 = _T_934 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1963 = _T_938 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1967 = _T_942 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1971 = _T_946 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1975 = _T_950 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1979 = _T_954 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1983 = _T_958 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1987 = _T_962 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1991 = _T_966 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1995 = _T_970 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1999 = _T_974 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2003 = _T_978 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2007 = _T_982 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2011 = _T_986 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2015 = _T_990 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2019 = _T_994 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2023 = _T_998 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2027 = _T_1002 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2031 = _T_1006 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2035 = _T_1010 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2039 = _T_1014 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2043 = _T_1018 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2047 = _T_1022 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2051 = _T_1026 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2055 = _T_1030 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2059 = _T_1034 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2063 = _T_1038 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2067 = _T_1042 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2071 = _T_1046 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2075 = _T_1050 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2079 = _T_1054 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2083 = _T_1058 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2087 = _T_1062 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2091 = _T_1066 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2095 = _T_1070 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2099 = _T_1074 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2103 = _T_1078 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2107 = _T_1082 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2111 = _T_1086 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2115 = _T_1090 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2119 = _T_1094 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2123 = _T_1098 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2127 = _T_1102 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2131 = _T_1106 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2135 = _T_1110 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2139 = _T_1114 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2143 = _T_1118 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2147 = _T_1122 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2151 = _T_1126 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2155 = _T_1130 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2159 = _T_1134 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2163 = _T_1138 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2167 = _T_1142 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2171 = _T_1146 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2175 = _T_1150 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2179 = _T_1154 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2183 = _T_1158 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2187 = _T_1162 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2191 = _T_1166 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2195 = _T_1170 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2199 = _T_1174 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2203 = _T_1178 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2207 = _T_1182 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2211 = _T_1186 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2215 = _T_1190 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2219 = _T_1194 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2223 = _T_1198 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2227 = _T_1202 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2231 = _T_1206 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2235 = _T_1210 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2239 = _T_1214 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2243 = _T_1218 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2247 = _T_1222 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2251 = _T_1226 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2255 = _T_1230 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2259 = _T_1234 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2263 = _T_1238 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2267 = _T_1242 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2271 = _T_1246 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2275 = _T_1250 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2279 = _T_1254 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2283 = _T_1258 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2287 = _T_1262 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2291 = _T_1266 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2295 = _T_1270 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2299 = _T_1274 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2303 = _T_1278 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2307 = _T_1282 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2311 = _T_1286 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2315 = _T_1290 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2319 = _T_1294 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2323 = _T_1298 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2327 = _T_1302 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2331 = _T_1306 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2335 = _T_1310 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2339 = _T_1314 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2343 = _T_1318 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2347 = _T_1322 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2351 = _T_1326 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2355 = _T_1330 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2359 = _T_1334 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2363 = _T_1338 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2367 = _T_1342 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2371 = _T_1346 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2375 = _T_1350 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2379 = _T_1354 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2383 = _T_1358 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2387 = _T_1362 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2391 = _T_1366 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2395 = _T_1370 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2399 = _T_1374 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2403 = _T_1378 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2407 = _T_1382 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2411 = _T_1386 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2415 = _T_1390 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2419 = _T_1394 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2423 = _T_1398 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2427 = _T_1402 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2431 = _T_1406 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2435 = _T_1410 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2439 = _T_1414 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2443 = _T_1418 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2447 = _T_1422 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2451 = _T_1426 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2455 = _T_1430 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2459 = _T_1434 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2463 = _T_1438 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2467 = _T_1442 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2471 = _T_1446 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2475 = _T_1450 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2479 = _T_1454 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2483 = _T_1458 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2487 = _T_1462 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2491 = _T_1466 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2495 = _T_1470 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2499 = _T_1474 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2503 = _T_1478 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2507 = _T_1482 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2511 = _T_1486 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2515 = _T_1490 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2519 = _T_1494 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2523 = _T_1498 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2527 = _T_1502 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2531 = _T_1506 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2535 = _T_1510 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2539 = _T_1514 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2543 = _T_1518 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2547 = _T_1522 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2551 = _T_1526 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2555 = _T_1530 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2559 = _T_1534 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2563 = _T_1538 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2567 = _T_1542 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2571 = _T_1546 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2575 = _T_1550 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2579 = _T_1554 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2583 = _T_1558 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2587 = _T_1562 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2591 = _T_1566 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2595 = _T_1570 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2599 = _T_1574 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2603 = _T_1578 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2607 = _T_1582 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2611 = _T_1586 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2615 = _T_1590 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2619 = _T_1594 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2623 = _T_1598 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2627 = _T_1602 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2631 = _T_1606 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2635 = _T_1610 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2639 = _T_1614 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2643 = _T_1618 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2647 = _T_1622 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2651 = _T_1626 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2655 = _T_1630 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2659 = _T_1634 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2663 = _T_1638 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2667 = _T_1642 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2671 = _T_1646 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2675 = _T_1650 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2679 = _T_1654 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2683 = _T_1658 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2687 = _T_1662 & _T_625; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_6788 = bht_wr_addr0[7:4] == 4'h0; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6790 = bht_wr_en0[0] & _T_6788; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6793 = bht_wr_addr2[7:4] == 4'h0; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6795 = bht_wr_en2[0] & _T_6793; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6799 = bht_wr_addr0[7:4] == 4'h1; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6801 = bht_wr_en0[0] & _T_6799; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6804 = bht_wr_addr2[7:4] == 4'h1; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6806 = bht_wr_en2[0] & _T_6804; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6810 = bht_wr_addr0[7:4] == 4'h2; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6812 = bht_wr_en0[0] & _T_6810; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6815 = bht_wr_addr2[7:4] == 4'h2; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6817 = bht_wr_en2[0] & _T_6815; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6821 = bht_wr_addr0[7:4] == 4'h3; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6823 = bht_wr_en0[0] & _T_6821; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6826 = bht_wr_addr2[7:4] == 4'h3; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6828 = bht_wr_en2[0] & _T_6826; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6832 = bht_wr_addr0[7:4] == 4'h4; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6834 = bht_wr_en0[0] & _T_6832; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6837 = bht_wr_addr2[7:4] == 4'h4; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6839 = bht_wr_en2[0] & _T_6837; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6843 = bht_wr_addr0[7:4] == 4'h5; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6845 = bht_wr_en0[0] & _T_6843; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6848 = bht_wr_addr2[7:4] == 4'h5; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6850 = bht_wr_en2[0] & _T_6848; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6854 = bht_wr_addr0[7:4] == 4'h6; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6856 = bht_wr_en0[0] & _T_6854; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6859 = bht_wr_addr2[7:4] == 4'h6; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6861 = bht_wr_en2[0] & _T_6859; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6865 = bht_wr_addr0[7:4] == 4'h7; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6867 = bht_wr_en0[0] & _T_6865; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6870 = bht_wr_addr2[7:4] == 4'h7; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6872 = bht_wr_en2[0] & _T_6870; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6876 = bht_wr_addr0[7:4] == 4'h8; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6878 = bht_wr_en0[0] & _T_6876; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6881 = bht_wr_addr2[7:4] == 4'h8; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6883 = bht_wr_en2[0] & _T_6881; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6887 = bht_wr_addr0[7:4] == 4'h9; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6889 = bht_wr_en0[0] & _T_6887; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6892 = bht_wr_addr2[7:4] == 4'h9; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6894 = bht_wr_en2[0] & _T_6892; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6898 = bht_wr_addr0[7:4] == 4'ha; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6900 = bht_wr_en0[0] & _T_6898; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6903 = bht_wr_addr2[7:4] == 4'ha; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6905 = bht_wr_en2[0] & _T_6903; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6909 = bht_wr_addr0[7:4] == 4'hb; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6911 = bht_wr_en0[0] & _T_6909; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6914 = bht_wr_addr2[7:4] == 4'hb; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6916 = bht_wr_en2[0] & _T_6914; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6920 = bht_wr_addr0[7:4] == 4'hc; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6922 = bht_wr_en0[0] & _T_6920; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6925 = bht_wr_addr2[7:4] == 4'hc; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6927 = bht_wr_en2[0] & _T_6925; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6931 = bht_wr_addr0[7:4] == 4'hd; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6933 = bht_wr_en0[0] & _T_6931; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6936 = bht_wr_addr2[7:4] == 4'hd; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6938 = bht_wr_en2[0] & _T_6936; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6942 = bht_wr_addr0[7:4] == 4'he; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6944 = bht_wr_en0[0] & _T_6942; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6947 = bht_wr_addr2[7:4] == 4'he; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6949 = bht_wr_en2[0] & _T_6947; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6953 = bht_wr_addr0[7:4] == 4'hf; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6955 = bht_wr_en0[0] & _T_6953; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6958 = bht_wr_addr2[7:4] == 4'hf; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6960 = bht_wr_en2[0] & _T_6958; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6966 = bht_wr_en0[1] & _T_6788; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6971 = bht_wr_en2[1] & _T_6793; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6977 = bht_wr_en0[1] & _T_6799; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6982 = bht_wr_en2[1] & _T_6804; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6988 = bht_wr_en0[1] & _T_6810; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6993 = bht_wr_en2[1] & _T_6815; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6999 = bht_wr_en0[1] & _T_6821; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7004 = bht_wr_en2[1] & _T_6826; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7010 = bht_wr_en0[1] & _T_6832; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7015 = bht_wr_en2[1] & _T_6837; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7021 = bht_wr_en0[1] & _T_6843; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7026 = bht_wr_en2[1] & _T_6848; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7032 = bht_wr_en0[1] & _T_6854; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7037 = bht_wr_en2[1] & _T_6859; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7043 = bht_wr_en0[1] & _T_6865; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7048 = bht_wr_en2[1] & _T_6870; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7054 = bht_wr_en0[1] & _T_6876; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7059 = bht_wr_en2[1] & _T_6881; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7065 = bht_wr_en0[1] & _T_6887; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7070 = bht_wr_en2[1] & _T_6892; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7076 = bht_wr_en0[1] & _T_6898; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7081 = bht_wr_en2[1] & _T_6903; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7087 = bht_wr_en0[1] & _T_6909; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7092 = bht_wr_en2[1] & _T_6914; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7098 = bht_wr_en0[1] & _T_6920; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7103 = bht_wr_en2[1] & _T_6925; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7109 = bht_wr_en0[1] & _T_6931; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7114 = bht_wr_en2[1] & _T_6936; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7120 = bht_wr_en0[1] & _T_6942; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7125 = bht_wr_en2[1] & _T_6947; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7131 = bht_wr_en0[1] & _T_6953; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_7136 = bht_wr_en2[1] & _T_6958; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_7140 = bht_wr_addr2[3:0] == 4'h0; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7141 = bht_wr_en2[0] & _T_7140; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7145 = _T_7141 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7149 = bht_wr_addr2[3:0] == 4'h1; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7150 = bht_wr_en2[0] & _T_7149; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7154 = _T_7150 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7158 = bht_wr_addr2[3:0] == 4'h2; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7159 = bht_wr_en2[0] & _T_7158; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7163 = _T_7159 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7167 = bht_wr_addr2[3:0] == 4'h3; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7168 = bht_wr_en2[0] & _T_7167; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7172 = _T_7168 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7176 = bht_wr_addr2[3:0] == 4'h4; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7177 = bht_wr_en2[0] & _T_7176; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7181 = _T_7177 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7185 = bht_wr_addr2[3:0] == 4'h5; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7186 = bht_wr_en2[0] & _T_7185; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7190 = _T_7186 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7194 = bht_wr_addr2[3:0] == 4'h6; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7195 = bht_wr_en2[0] & _T_7194; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7199 = _T_7195 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7203 = bht_wr_addr2[3:0] == 4'h7; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7204 = bht_wr_en2[0] & _T_7203; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7208 = _T_7204 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7212 = bht_wr_addr2[3:0] == 4'h8; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7213 = bht_wr_en2[0] & _T_7212; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7217 = _T_7213 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7221 = bht_wr_addr2[3:0] == 4'h9; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7222 = bht_wr_en2[0] & _T_7221; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7226 = _T_7222 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7230 = bht_wr_addr2[3:0] == 4'ha; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7231 = bht_wr_en2[0] & _T_7230; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7235 = _T_7231 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7239 = bht_wr_addr2[3:0] == 4'hb; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7240 = bht_wr_en2[0] & _T_7239; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7244 = _T_7240 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7248 = bht_wr_addr2[3:0] == 4'hc; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7249 = bht_wr_en2[0] & _T_7248; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7253 = _T_7249 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7257 = bht_wr_addr2[3:0] == 4'hd; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7258 = bht_wr_en2[0] & _T_7257; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7262 = _T_7258 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7266 = bht_wr_addr2[3:0] == 4'he; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7267 = bht_wr_en2[0] & _T_7266; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7271 = _T_7267 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7275 = bht_wr_addr2[3:0] == 4'hf; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_7276 = bht_wr_en2[0] & _T_7275; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_7280 = _T_7276 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7289 = _T_7141 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7298 = _T_7150 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7307 = _T_7159 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7316 = _T_7168 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7325 = _T_7177 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7334 = _T_7186 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7343 = _T_7195 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7352 = _T_7204 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7361 = _T_7213 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7370 = _T_7222 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7379 = _T_7231 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7388 = _T_7240 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7397 = _T_7249 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7406 = _T_7258 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7415 = _T_7267 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7424 = _T_7276 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7433 = _T_7141 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7442 = _T_7150 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7451 = _T_7159 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7460 = _T_7168 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7469 = _T_7177 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7478 = _T_7186 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7487 = _T_7195 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7496 = _T_7204 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7505 = _T_7213 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7514 = _T_7222 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7523 = _T_7231 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7532 = _T_7240 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7541 = _T_7249 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7550 = _T_7258 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7559 = _T_7267 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7568 = _T_7276 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7577 = _T_7141 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7586 = _T_7150 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7595 = _T_7159 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7604 = _T_7168 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7613 = _T_7177 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7622 = _T_7186 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7631 = _T_7195 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7640 = _T_7204 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7649 = _T_7213 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7658 = _T_7222 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7667 = _T_7231 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7676 = _T_7240 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7685 = _T_7249 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7694 = _T_7258 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7703 = _T_7267 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7712 = _T_7276 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7721 = _T_7141 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7730 = _T_7150 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7739 = _T_7159 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7748 = _T_7168 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7757 = _T_7177 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7766 = _T_7186 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7775 = _T_7195 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7784 = _T_7204 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7793 = _T_7213 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7802 = _T_7222 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7811 = _T_7231 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7820 = _T_7240 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7829 = _T_7249 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7838 = _T_7258 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7847 = _T_7267 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7856 = _T_7276 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7865 = _T_7141 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7874 = _T_7150 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7883 = _T_7159 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7892 = _T_7168 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7901 = _T_7177 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7910 = _T_7186 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7919 = _T_7195 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7928 = _T_7204 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7937 = _T_7213 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7946 = _T_7222 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7955 = _T_7231 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7964 = _T_7240 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7973 = _T_7249 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7982 = _T_7258 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7991 = _T_7267 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8000 = _T_7276 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8009 = _T_7141 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8018 = _T_7150 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8027 = _T_7159 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8036 = _T_7168 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8045 = _T_7177 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8054 = _T_7186 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8063 = _T_7195 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8072 = _T_7204 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8081 = _T_7213 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8090 = _T_7222 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8099 = _T_7231 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8108 = _T_7240 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8117 = _T_7249 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8126 = _T_7258 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8135 = _T_7267 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8144 = _T_7276 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8153 = _T_7141 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8162 = _T_7150 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8171 = _T_7159 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8180 = _T_7168 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8189 = _T_7177 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8198 = _T_7186 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8207 = _T_7195 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8216 = _T_7204 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8225 = _T_7213 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8234 = _T_7222 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8243 = _T_7231 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8252 = _T_7240 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8261 = _T_7249 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8270 = _T_7258 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8279 = _T_7267 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8288 = _T_7276 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8297 = _T_7141 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8306 = _T_7150 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8315 = _T_7159 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8324 = _T_7168 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8333 = _T_7177 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8342 = _T_7186 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8351 = _T_7195 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8360 = _T_7204 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8369 = _T_7213 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8378 = _T_7222 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8387 = _T_7231 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8396 = _T_7240 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8405 = _T_7249 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8414 = _T_7258 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8423 = _T_7267 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8432 = _T_7276 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8441 = _T_7141 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8450 = _T_7150 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8459 = _T_7159 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8468 = _T_7168 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8477 = _T_7177 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8486 = _T_7186 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8495 = _T_7195 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8504 = _T_7204 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8513 = _T_7213 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8522 = _T_7222 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8531 = _T_7231 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8540 = _T_7240 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8549 = _T_7249 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8558 = _T_7258 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8567 = _T_7267 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8576 = _T_7276 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8585 = _T_7141 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8594 = _T_7150 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8603 = _T_7159 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8612 = _T_7168 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8621 = _T_7177 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8630 = _T_7186 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8639 = _T_7195 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8648 = _T_7204 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8657 = _T_7213 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8666 = _T_7222 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8675 = _T_7231 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8684 = _T_7240 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8693 = _T_7249 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8702 = _T_7258 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8711 = _T_7267 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8720 = _T_7276 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8729 = _T_7141 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8738 = _T_7150 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8747 = _T_7159 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8756 = _T_7168 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8765 = _T_7177 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8774 = _T_7186 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8783 = _T_7195 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8792 = _T_7204 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8801 = _T_7213 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8810 = _T_7222 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8819 = _T_7231 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8828 = _T_7240 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8837 = _T_7249 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8846 = _T_7258 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8855 = _T_7267 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8864 = _T_7276 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8873 = _T_7141 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8882 = _T_7150 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8891 = _T_7159 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8900 = _T_7168 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8909 = _T_7177 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8918 = _T_7186 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8927 = _T_7195 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8936 = _T_7204 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8945 = _T_7213 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8954 = _T_7222 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8963 = _T_7231 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8972 = _T_7240 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8981 = _T_7249 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8990 = _T_7258 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8999 = _T_7267 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9008 = _T_7276 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9017 = _T_7141 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9026 = _T_7150 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9035 = _T_7159 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9044 = _T_7168 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9053 = _T_7177 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9062 = _T_7186 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9071 = _T_7195 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9080 = _T_7204 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9089 = _T_7213 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9098 = _T_7222 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9107 = _T_7231 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9116 = _T_7240 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9125 = _T_7249 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9134 = _T_7258 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9143 = _T_7267 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9152 = _T_7276 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9161 = _T_7141 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9170 = _T_7150 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9179 = _T_7159 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9188 = _T_7168 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9197 = _T_7177 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9206 = _T_7186 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9215 = _T_7195 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9224 = _T_7204 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9233 = _T_7213 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9242 = _T_7222 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9251 = _T_7231 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9260 = _T_7240 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9269 = _T_7249 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9278 = _T_7258 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9287 = _T_7267 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9296 = _T_7276 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9305 = _T_7141 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9314 = _T_7150 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9323 = _T_7159 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9332 = _T_7168 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9341 = _T_7177 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9350 = _T_7186 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9359 = _T_7195 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9368 = _T_7204 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9377 = _T_7213 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9386 = _T_7222 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9395 = _T_7231 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9404 = _T_7240 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9413 = _T_7249 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9422 = _T_7258 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9431 = _T_7267 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9440 = _T_7276 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9445 = bht_wr_en2[1] & _T_7140; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9449 = _T_9445 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9454 = bht_wr_en2[1] & _T_7149; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9458 = _T_9454 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9463 = bht_wr_en2[1] & _T_7158; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9467 = _T_9463 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9472 = bht_wr_en2[1] & _T_7167; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9476 = _T_9472 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9481 = bht_wr_en2[1] & _T_7176; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9485 = _T_9481 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9490 = bht_wr_en2[1] & _T_7185; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9494 = _T_9490 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9499 = bht_wr_en2[1] & _T_7194; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9503 = _T_9499 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9508 = bht_wr_en2[1] & _T_7203; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9512 = _T_9508 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9517 = bht_wr_en2[1] & _T_7212; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9521 = _T_9517 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9526 = bht_wr_en2[1] & _T_7221; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9530 = _T_9526 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9535 = bht_wr_en2[1] & _T_7230; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9539 = _T_9535 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9544 = bht_wr_en2[1] & _T_7239; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9548 = _T_9544 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9553 = bht_wr_en2[1] & _T_7248; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9557 = _T_9553 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9562 = bht_wr_en2[1] & _T_7257; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9566 = _T_9562 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9571 = bht_wr_en2[1] & _T_7266; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9575 = _T_9571 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9580 = bht_wr_en2[1] & _T_7275; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9584 = _T_9580 & _T_6793; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9593 = _T_9445 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9602 = _T_9454 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9611 = _T_9463 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9620 = _T_9472 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9629 = _T_9481 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9638 = _T_9490 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9647 = _T_9499 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9656 = _T_9508 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9665 = _T_9517 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9674 = _T_9526 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9683 = _T_9535 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9692 = _T_9544 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9701 = _T_9553 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9710 = _T_9562 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9719 = _T_9571 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9728 = _T_9580 & _T_6804; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9737 = _T_9445 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9746 = _T_9454 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9755 = _T_9463 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9764 = _T_9472 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9773 = _T_9481 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9782 = _T_9490 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9791 = _T_9499 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9800 = _T_9508 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9809 = _T_9517 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9818 = _T_9526 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9827 = _T_9535 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9836 = _T_9544 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9845 = _T_9553 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9854 = _T_9562 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9863 = _T_9571 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9872 = _T_9580 & _T_6815; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9881 = _T_9445 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9890 = _T_9454 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9899 = _T_9463 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9908 = _T_9472 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9917 = _T_9481 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9926 = _T_9490 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9935 = _T_9499 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9944 = _T_9508 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9953 = _T_9517 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9962 = _T_9526 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9971 = _T_9535 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9980 = _T_9544 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9989 = _T_9553 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9998 = _T_9562 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10007 = _T_9571 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10016 = _T_9580 & _T_6826; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10025 = _T_9445 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10034 = _T_9454 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10043 = _T_9463 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10052 = _T_9472 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10061 = _T_9481 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10070 = _T_9490 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10079 = _T_9499 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10088 = _T_9508 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10097 = _T_9517 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10106 = _T_9526 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10115 = _T_9535 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10124 = _T_9544 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10133 = _T_9553 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10142 = _T_9562 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10151 = _T_9571 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10160 = _T_9580 & _T_6837; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10169 = _T_9445 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10178 = _T_9454 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10187 = _T_9463 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10196 = _T_9472 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10205 = _T_9481 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10214 = _T_9490 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10223 = _T_9499 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10232 = _T_9508 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10241 = _T_9517 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10250 = _T_9526 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10259 = _T_9535 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10268 = _T_9544 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10277 = _T_9553 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10286 = _T_9562 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10295 = _T_9571 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10304 = _T_9580 & _T_6848; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10313 = _T_9445 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10322 = _T_9454 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10331 = _T_9463 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10340 = _T_9472 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10349 = _T_9481 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10358 = _T_9490 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10367 = _T_9499 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10376 = _T_9508 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10385 = _T_9517 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10394 = _T_9526 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10403 = _T_9535 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10412 = _T_9544 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10421 = _T_9553 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10430 = _T_9562 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10439 = _T_9571 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10448 = _T_9580 & _T_6859; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10457 = _T_9445 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10466 = _T_9454 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10475 = _T_9463 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10484 = _T_9472 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10493 = _T_9481 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10502 = _T_9490 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10511 = _T_9499 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10520 = _T_9508 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10529 = _T_9517 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10538 = _T_9526 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10547 = _T_9535 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10556 = _T_9544 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10565 = _T_9553 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10574 = _T_9562 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10583 = _T_9571 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10592 = _T_9580 & _T_6870; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10601 = _T_9445 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10610 = _T_9454 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10619 = _T_9463 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10628 = _T_9472 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10637 = _T_9481 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10646 = _T_9490 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10655 = _T_9499 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10664 = _T_9508 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10673 = _T_9517 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10682 = _T_9526 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10691 = _T_9535 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10700 = _T_9544 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10709 = _T_9553 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10718 = _T_9562 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10727 = _T_9571 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10736 = _T_9580 & _T_6881; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10745 = _T_9445 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10754 = _T_9454 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10763 = _T_9463 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10772 = _T_9472 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10781 = _T_9481 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10790 = _T_9490 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10799 = _T_9499 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10808 = _T_9508 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10817 = _T_9517 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10826 = _T_9526 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10835 = _T_9535 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10844 = _T_9544 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10853 = _T_9553 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10862 = _T_9562 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10871 = _T_9571 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10880 = _T_9580 & _T_6892; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10889 = _T_9445 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10898 = _T_9454 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10907 = _T_9463 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10916 = _T_9472 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10925 = _T_9481 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10934 = _T_9490 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10943 = _T_9499 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10952 = _T_9508 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10961 = _T_9517 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10970 = _T_9526 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10979 = _T_9535 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10988 = _T_9544 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10997 = _T_9553 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11006 = _T_9562 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11015 = _T_9571 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11024 = _T_9580 & _T_6903; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11033 = _T_9445 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11042 = _T_9454 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11051 = _T_9463 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11060 = _T_9472 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11069 = _T_9481 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11078 = _T_9490 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11087 = _T_9499 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11096 = _T_9508 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11105 = _T_9517 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11114 = _T_9526 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11123 = _T_9535 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11132 = _T_9544 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11141 = _T_9553 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11150 = _T_9562 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11159 = _T_9571 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11168 = _T_9580 & _T_6914; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11177 = _T_9445 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11186 = _T_9454 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11195 = _T_9463 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11204 = _T_9472 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11213 = _T_9481 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11222 = _T_9490 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11231 = _T_9499 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11240 = _T_9508 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11249 = _T_9517 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11258 = _T_9526 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11267 = _T_9535 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11276 = _T_9544 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11285 = _T_9553 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11294 = _T_9562 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11303 = _T_9571 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11312 = _T_9580 & _T_6925; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11321 = _T_9445 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11330 = _T_9454 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11339 = _T_9463 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11348 = _T_9472 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11357 = _T_9481 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11366 = _T_9490 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11375 = _T_9499 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11384 = _T_9508 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11393 = _T_9517 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11402 = _T_9526 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11411 = _T_9535 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11420 = _T_9544 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11429 = _T_9553 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11438 = _T_9562 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11447 = _T_9571 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11456 = _T_9580 & _T_6936; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11465 = _T_9445 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11474 = _T_9454 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11483 = _T_9463 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11492 = _T_9472 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11501 = _T_9481 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11510 = _T_9490 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11519 = _T_9499 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11528 = _T_9508 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11537 = _T_9517 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11546 = _T_9526 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11555 = _T_9535 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11564 = _T_9544 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11573 = _T_9553 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11582 = _T_9562 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11591 = _T_9571 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11600 = _T_9580 & _T_6947; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11609 = _T_9445 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11618 = _T_9454 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11627 = _T_9463 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11636 = _T_9472 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11645 = _T_9481 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11654 = _T_9490 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11663 = _T_9499 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11672 = _T_9508 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11681 = _T_9517 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11690 = _T_9526 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11699 = _T_9535 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11708 = _T_9544 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11717 = _T_9553 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11726 = _T_9562 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11735 = _T_9571 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11744 = _T_9580 & _T_6958; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11748 = bht_wr_addr0[3:0] == 4'h0; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11749 = bht_wr_en0[0] & _T_11748; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11753 = _T_11749 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_0 = _T_11753 | _T_7145; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11765 = bht_wr_addr0[3:0] == 4'h1; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11766 = bht_wr_en0[0] & _T_11765; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11770 = _T_11766 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_1 = _T_11770 | _T_7154; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11782 = bht_wr_addr0[3:0] == 4'h2; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11783 = bht_wr_en0[0] & _T_11782; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11787 = _T_11783 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_2 = _T_11787 | _T_7163; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11799 = bht_wr_addr0[3:0] == 4'h3; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11800 = bht_wr_en0[0] & _T_11799; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11804 = _T_11800 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_3 = _T_11804 | _T_7172; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11816 = bht_wr_addr0[3:0] == 4'h4; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11817 = bht_wr_en0[0] & _T_11816; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11821 = _T_11817 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_4 = _T_11821 | _T_7181; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11833 = bht_wr_addr0[3:0] == 4'h5; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11834 = bht_wr_en0[0] & _T_11833; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11838 = _T_11834 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_5 = _T_11838 | _T_7190; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11850 = bht_wr_addr0[3:0] == 4'h6; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11851 = bht_wr_en0[0] & _T_11850; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11855 = _T_11851 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_6 = _T_11855 | _T_7199; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11867 = bht_wr_addr0[3:0] == 4'h7; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11868 = bht_wr_en0[0] & _T_11867; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11872 = _T_11868 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_7 = _T_11872 | _T_7208; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11884 = bht_wr_addr0[3:0] == 4'h8; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11885 = bht_wr_en0[0] & _T_11884; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11889 = _T_11885 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_8 = _T_11889 | _T_7217; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11901 = bht_wr_addr0[3:0] == 4'h9; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11902 = bht_wr_en0[0] & _T_11901; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11906 = _T_11902 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_9 = _T_11906 | _T_7226; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11918 = bht_wr_addr0[3:0] == 4'ha; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11919 = bht_wr_en0[0] & _T_11918; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11923 = _T_11919 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_10 = _T_11923 | _T_7235; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11935 = bht_wr_addr0[3:0] == 4'hb; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11936 = bht_wr_en0[0] & _T_11935; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11940 = _T_11936 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_11 = _T_11940 | _T_7244; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11952 = bht_wr_addr0[3:0] == 4'hc; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11953 = bht_wr_en0[0] & _T_11952; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11957 = _T_11953 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_12 = _T_11957 | _T_7253; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11969 = bht_wr_addr0[3:0] == 4'hd; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11970 = bht_wr_en0[0] & _T_11969; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11974 = _T_11970 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_13 = _T_11974 | _T_7262; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11986 = bht_wr_addr0[3:0] == 4'he; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11987 = bht_wr_en0[0] & _T_11986; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11991 = _T_11987 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_14 = _T_11991 | _T_7271; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12003 = bht_wr_addr0[3:0] == 4'hf; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_12004 = bht_wr_en0[0] & _T_12003; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_12008 = _T_12004 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_15 = _T_12008 | _T_7280; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12025 = _T_11749 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_0 = _T_12025 | _T_7289; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12042 = _T_11766 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_1 = _T_12042 | _T_7298; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12059 = _T_11783 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_2 = _T_12059 | _T_7307; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12076 = _T_11800 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_3 = _T_12076 | _T_7316; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12093 = _T_11817 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_4 = _T_12093 | _T_7325; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12110 = _T_11834 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_5 = _T_12110 | _T_7334; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12127 = _T_11851 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_6 = _T_12127 | _T_7343; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12144 = _T_11868 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_7 = _T_12144 | _T_7352; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12161 = _T_11885 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_8 = _T_12161 | _T_7361; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12178 = _T_11902 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_9 = _T_12178 | _T_7370; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12195 = _T_11919 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_10 = _T_12195 | _T_7379; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12212 = _T_11936 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_11 = _T_12212 | _T_7388; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12229 = _T_11953 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_12 = _T_12229 | _T_7397; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12246 = _T_11970 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_13 = _T_12246 | _T_7406; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12263 = _T_11987 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_14 = _T_12263 | _T_7415; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12280 = _T_12004 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_15 = _T_12280 | _T_7424; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12297 = _T_11749 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_0 = _T_12297 | _T_7433; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12314 = _T_11766 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_1 = _T_12314 | _T_7442; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12331 = _T_11783 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_2 = _T_12331 | _T_7451; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12348 = _T_11800 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_3 = _T_12348 | _T_7460; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12365 = _T_11817 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_4 = _T_12365 | _T_7469; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12382 = _T_11834 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_5 = _T_12382 | _T_7478; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12399 = _T_11851 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_6 = _T_12399 | _T_7487; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12416 = _T_11868 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_7 = _T_12416 | _T_7496; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12433 = _T_11885 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_8 = _T_12433 | _T_7505; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12450 = _T_11902 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_9 = _T_12450 | _T_7514; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12467 = _T_11919 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_10 = _T_12467 | _T_7523; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12484 = _T_11936 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_11 = _T_12484 | _T_7532; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12501 = _T_11953 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_12 = _T_12501 | _T_7541; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12518 = _T_11970 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_13 = _T_12518 | _T_7550; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12535 = _T_11987 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_14 = _T_12535 | _T_7559; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12552 = _T_12004 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_15 = _T_12552 | _T_7568; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12569 = _T_11749 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_0 = _T_12569 | _T_7577; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12586 = _T_11766 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_1 = _T_12586 | _T_7586; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12603 = _T_11783 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_2 = _T_12603 | _T_7595; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12620 = _T_11800 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_3 = _T_12620 | _T_7604; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12637 = _T_11817 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_4 = _T_12637 | _T_7613; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12654 = _T_11834 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_5 = _T_12654 | _T_7622; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12671 = _T_11851 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_6 = _T_12671 | _T_7631; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12688 = _T_11868 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_7 = _T_12688 | _T_7640; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12705 = _T_11885 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_8 = _T_12705 | _T_7649; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12722 = _T_11902 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_9 = _T_12722 | _T_7658; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12739 = _T_11919 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_10 = _T_12739 | _T_7667; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12756 = _T_11936 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_11 = _T_12756 | _T_7676; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12773 = _T_11953 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_12 = _T_12773 | _T_7685; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12790 = _T_11970 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_13 = _T_12790 | _T_7694; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12807 = _T_11987 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_14 = _T_12807 | _T_7703; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12824 = _T_12004 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_15 = _T_12824 | _T_7712; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12841 = _T_11749 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_0 = _T_12841 | _T_7721; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12858 = _T_11766 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_1 = _T_12858 | _T_7730; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12875 = _T_11783 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_2 = _T_12875 | _T_7739; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12892 = _T_11800 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_3 = _T_12892 | _T_7748; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12909 = _T_11817 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_4 = _T_12909 | _T_7757; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12926 = _T_11834 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_5 = _T_12926 | _T_7766; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12943 = _T_11851 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_6 = _T_12943 | _T_7775; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12960 = _T_11868 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_7 = _T_12960 | _T_7784; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12977 = _T_11885 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_8 = _T_12977 | _T_7793; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12994 = _T_11902 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_9 = _T_12994 | _T_7802; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13011 = _T_11919 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_10 = _T_13011 | _T_7811; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13028 = _T_11936 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_11 = _T_13028 | _T_7820; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13045 = _T_11953 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_12 = _T_13045 | _T_7829; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13062 = _T_11970 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_13 = _T_13062 | _T_7838; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13079 = _T_11987 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_14 = _T_13079 | _T_7847; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13096 = _T_12004 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_15 = _T_13096 | _T_7856; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13113 = _T_11749 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_0 = _T_13113 | _T_7865; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13130 = _T_11766 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_1 = _T_13130 | _T_7874; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13147 = _T_11783 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_2 = _T_13147 | _T_7883; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13164 = _T_11800 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_3 = _T_13164 | _T_7892; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13181 = _T_11817 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_4 = _T_13181 | _T_7901; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13198 = _T_11834 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_5 = _T_13198 | _T_7910; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13215 = _T_11851 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_6 = _T_13215 | _T_7919; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13232 = _T_11868 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_7 = _T_13232 | _T_7928; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13249 = _T_11885 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_8 = _T_13249 | _T_7937; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13266 = _T_11902 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_9 = _T_13266 | _T_7946; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13283 = _T_11919 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_10 = _T_13283 | _T_7955; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13300 = _T_11936 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_11 = _T_13300 | _T_7964; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13317 = _T_11953 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_12 = _T_13317 | _T_7973; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13334 = _T_11970 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_13 = _T_13334 | _T_7982; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13351 = _T_11987 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_14 = _T_13351 | _T_7991; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13368 = _T_12004 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_15 = _T_13368 | _T_8000; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13385 = _T_11749 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_0 = _T_13385 | _T_8009; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13402 = _T_11766 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_1 = _T_13402 | _T_8018; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13419 = _T_11783 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_2 = _T_13419 | _T_8027; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13436 = _T_11800 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_3 = _T_13436 | _T_8036; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13453 = _T_11817 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_4 = _T_13453 | _T_8045; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13470 = _T_11834 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_5 = _T_13470 | _T_8054; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13487 = _T_11851 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_6 = _T_13487 | _T_8063; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13504 = _T_11868 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_7 = _T_13504 | _T_8072; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13521 = _T_11885 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_8 = _T_13521 | _T_8081; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13538 = _T_11902 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_9 = _T_13538 | _T_8090; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13555 = _T_11919 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_10 = _T_13555 | _T_8099; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13572 = _T_11936 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_11 = _T_13572 | _T_8108; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13589 = _T_11953 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_12 = _T_13589 | _T_8117; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13606 = _T_11970 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_13 = _T_13606 | _T_8126; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13623 = _T_11987 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_14 = _T_13623 | _T_8135; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13640 = _T_12004 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_15 = _T_13640 | _T_8144; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13657 = _T_11749 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_0 = _T_13657 | _T_8153; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13674 = _T_11766 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_1 = _T_13674 | _T_8162; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13691 = _T_11783 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_2 = _T_13691 | _T_8171; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13708 = _T_11800 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_3 = _T_13708 | _T_8180; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13725 = _T_11817 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_4 = _T_13725 | _T_8189; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13742 = _T_11834 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_5 = _T_13742 | _T_8198; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13759 = _T_11851 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_6 = _T_13759 | _T_8207; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13776 = _T_11868 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_7 = _T_13776 | _T_8216; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13793 = _T_11885 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_8 = _T_13793 | _T_8225; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13810 = _T_11902 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_9 = _T_13810 | _T_8234; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13827 = _T_11919 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_10 = _T_13827 | _T_8243; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13844 = _T_11936 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_11 = _T_13844 | _T_8252; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13861 = _T_11953 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_12 = _T_13861 | _T_8261; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13878 = _T_11970 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_13 = _T_13878 | _T_8270; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13895 = _T_11987 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_14 = _T_13895 | _T_8279; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13912 = _T_12004 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_15 = _T_13912 | _T_8288; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13929 = _T_11749 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_0 = _T_13929 | _T_8297; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13946 = _T_11766 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_1 = _T_13946 | _T_8306; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13963 = _T_11783 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_2 = _T_13963 | _T_8315; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13980 = _T_11800 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_3 = _T_13980 | _T_8324; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13997 = _T_11817 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_4 = _T_13997 | _T_8333; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14014 = _T_11834 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_5 = _T_14014 | _T_8342; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14031 = _T_11851 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_6 = _T_14031 | _T_8351; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14048 = _T_11868 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_7 = _T_14048 | _T_8360; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14065 = _T_11885 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_8 = _T_14065 | _T_8369; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14082 = _T_11902 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_9 = _T_14082 | _T_8378; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14099 = _T_11919 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_10 = _T_14099 | _T_8387; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14116 = _T_11936 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_11 = _T_14116 | _T_8396; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14133 = _T_11953 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_12 = _T_14133 | _T_8405; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14150 = _T_11970 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_13 = _T_14150 | _T_8414; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14167 = _T_11987 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_14 = _T_14167 | _T_8423; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14184 = _T_12004 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_15 = _T_14184 | _T_8432; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14201 = _T_11749 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_0 = _T_14201 | _T_8441; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14218 = _T_11766 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_1 = _T_14218 | _T_8450; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14235 = _T_11783 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_2 = _T_14235 | _T_8459; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14252 = _T_11800 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_3 = _T_14252 | _T_8468; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14269 = _T_11817 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_4 = _T_14269 | _T_8477; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14286 = _T_11834 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_5 = _T_14286 | _T_8486; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14303 = _T_11851 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_6 = _T_14303 | _T_8495; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14320 = _T_11868 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_7 = _T_14320 | _T_8504; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14337 = _T_11885 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_8 = _T_14337 | _T_8513; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14354 = _T_11902 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_9 = _T_14354 | _T_8522; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14371 = _T_11919 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_10 = _T_14371 | _T_8531; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14388 = _T_11936 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_11 = _T_14388 | _T_8540; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14405 = _T_11953 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_12 = _T_14405 | _T_8549; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14422 = _T_11970 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_13 = _T_14422 | _T_8558; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14439 = _T_11987 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_14 = _T_14439 | _T_8567; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14456 = _T_12004 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_15 = _T_14456 | _T_8576; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14473 = _T_11749 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_0 = _T_14473 | _T_8585; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14490 = _T_11766 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_1 = _T_14490 | _T_8594; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14507 = _T_11783 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_2 = _T_14507 | _T_8603; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14524 = _T_11800 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_3 = _T_14524 | _T_8612; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14541 = _T_11817 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_4 = _T_14541 | _T_8621; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14558 = _T_11834 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_5 = _T_14558 | _T_8630; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14575 = _T_11851 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_6 = _T_14575 | _T_8639; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14592 = _T_11868 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_7 = _T_14592 | _T_8648; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14609 = _T_11885 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_8 = _T_14609 | _T_8657; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14626 = _T_11902 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_9 = _T_14626 | _T_8666; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14643 = _T_11919 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_10 = _T_14643 | _T_8675; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14660 = _T_11936 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_11 = _T_14660 | _T_8684; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14677 = _T_11953 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_12 = _T_14677 | _T_8693; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14694 = _T_11970 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_13 = _T_14694 | _T_8702; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14711 = _T_11987 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_14 = _T_14711 | _T_8711; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14728 = _T_12004 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_15 = _T_14728 | _T_8720; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14745 = _T_11749 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_0 = _T_14745 | _T_8729; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14762 = _T_11766 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_1 = _T_14762 | _T_8738; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14779 = _T_11783 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_2 = _T_14779 | _T_8747; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14796 = _T_11800 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_3 = _T_14796 | _T_8756; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14813 = _T_11817 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_4 = _T_14813 | _T_8765; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14830 = _T_11834 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_5 = _T_14830 | _T_8774; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14847 = _T_11851 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_6 = _T_14847 | _T_8783; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14864 = _T_11868 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_7 = _T_14864 | _T_8792; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14881 = _T_11885 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_8 = _T_14881 | _T_8801; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14898 = _T_11902 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_9 = _T_14898 | _T_8810; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14915 = _T_11919 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_10 = _T_14915 | _T_8819; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14932 = _T_11936 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_11 = _T_14932 | _T_8828; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14949 = _T_11953 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_12 = _T_14949 | _T_8837; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14966 = _T_11970 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_13 = _T_14966 | _T_8846; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14983 = _T_11987 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_14 = _T_14983 | _T_8855; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15000 = _T_12004 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_15 = _T_15000 | _T_8864; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15017 = _T_11749 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_0 = _T_15017 | _T_8873; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15034 = _T_11766 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_1 = _T_15034 | _T_8882; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15051 = _T_11783 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_2 = _T_15051 | _T_8891; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15068 = _T_11800 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_3 = _T_15068 | _T_8900; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15085 = _T_11817 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_4 = _T_15085 | _T_8909; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15102 = _T_11834 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_5 = _T_15102 | _T_8918; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15119 = _T_11851 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_6 = _T_15119 | _T_8927; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15136 = _T_11868 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_7 = _T_15136 | _T_8936; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15153 = _T_11885 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_8 = _T_15153 | _T_8945; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15170 = _T_11902 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_9 = _T_15170 | _T_8954; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15187 = _T_11919 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_10 = _T_15187 | _T_8963; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15204 = _T_11936 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_11 = _T_15204 | _T_8972; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15221 = _T_11953 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_12 = _T_15221 | _T_8981; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15238 = _T_11970 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_13 = _T_15238 | _T_8990; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15255 = _T_11987 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_14 = _T_15255 | _T_8999; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15272 = _T_12004 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_15 = _T_15272 | _T_9008; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15289 = _T_11749 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_0 = _T_15289 | _T_9017; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15306 = _T_11766 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_1 = _T_15306 | _T_9026; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15323 = _T_11783 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_2 = _T_15323 | _T_9035; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15340 = _T_11800 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_3 = _T_15340 | _T_9044; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15357 = _T_11817 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_4 = _T_15357 | _T_9053; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15374 = _T_11834 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_5 = _T_15374 | _T_9062; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15391 = _T_11851 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_6 = _T_15391 | _T_9071; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15408 = _T_11868 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_7 = _T_15408 | _T_9080; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15425 = _T_11885 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_8 = _T_15425 | _T_9089; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15442 = _T_11902 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_9 = _T_15442 | _T_9098; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15459 = _T_11919 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_10 = _T_15459 | _T_9107; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15476 = _T_11936 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_11 = _T_15476 | _T_9116; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15493 = _T_11953 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_12 = _T_15493 | _T_9125; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15510 = _T_11970 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_13 = _T_15510 | _T_9134; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15527 = _T_11987 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_14 = _T_15527 | _T_9143; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15544 = _T_12004 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_15 = _T_15544 | _T_9152; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15561 = _T_11749 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_0 = _T_15561 | _T_9161; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15578 = _T_11766 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_1 = _T_15578 | _T_9170; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15595 = _T_11783 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_2 = _T_15595 | _T_9179; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15612 = _T_11800 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_3 = _T_15612 | _T_9188; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15629 = _T_11817 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_4 = _T_15629 | _T_9197; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15646 = _T_11834 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_5 = _T_15646 | _T_9206; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15663 = _T_11851 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_6 = _T_15663 | _T_9215; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15680 = _T_11868 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_7 = _T_15680 | _T_9224; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15697 = _T_11885 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_8 = _T_15697 | _T_9233; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15714 = _T_11902 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_9 = _T_15714 | _T_9242; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15731 = _T_11919 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_10 = _T_15731 | _T_9251; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15748 = _T_11936 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_11 = _T_15748 | _T_9260; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15765 = _T_11953 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_12 = _T_15765 | _T_9269; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15782 = _T_11970 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_13 = _T_15782 | _T_9278; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15799 = _T_11987 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_14 = _T_15799 | _T_9287; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15816 = _T_12004 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_15 = _T_15816 | _T_9296; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15833 = _T_11749 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_0 = _T_15833 | _T_9305; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15850 = _T_11766 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_1 = _T_15850 | _T_9314; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15867 = _T_11783 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_2 = _T_15867 | _T_9323; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15884 = _T_11800 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_3 = _T_15884 | _T_9332; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15901 = _T_11817 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_4 = _T_15901 | _T_9341; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15918 = _T_11834 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_5 = _T_15918 | _T_9350; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15935 = _T_11851 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_6 = _T_15935 | _T_9359; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15952 = _T_11868 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_7 = _T_15952 | _T_9368; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15969 = _T_11885 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_8 = _T_15969 | _T_9377; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15986 = _T_11902 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_9 = _T_15986 | _T_9386; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16003 = _T_11919 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_10 = _T_16003 | _T_9395; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16020 = _T_11936 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_11 = _T_16020 | _T_9404; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16037 = _T_11953 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_12 = _T_16037 | _T_9413; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16054 = _T_11970 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_13 = _T_16054 | _T_9422; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16071 = _T_11987 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_14 = _T_16071 | _T_9431; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16088 = _T_12004 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_15 = _T_16088 | _T_9440; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16101 = bht_wr_en0[1] & _T_11748; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16105 = _T_16101 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_0 = _T_16105 | _T_9449; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16118 = bht_wr_en0[1] & _T_11765; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16122 = _T_16118 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_1 = _T_16122 | _T_9458; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16135 = bht_wr_en0[1] & _T_11782; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16139 = _T_16135 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_2 = _T_16139 | _T_9467; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16152 = bht_wr_en0[1] & _T_11799; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16156 = _T_16152 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_3 = _T_16156 | _T_9476; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16169 = bht_wr_en0[1] & _T_11816; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16173 = _T_16169 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_4 = _T_16173 | _T_9485; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16186 = bht_wr_en0[1] & _T_11833; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16190 = _T_16186 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_5 = _T_16190 | _T_9494; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16203 = bht_wr_en0[1] & _T_11850; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16207 = _T_16203 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_6 = _T_16207 | _T_9503; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16220 = bht_wr_en0[1] & _T_11867; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16224 = _T_16220 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_7 = _T_16224 | _T_9512; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16237 = bht_wr_en0[1] & _T_11884; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16241 = _T_16237 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_8 = _T_16241 | _T_9521; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16254 = bht_wr_en0[1] & _T_11901; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16258 = _T_16254 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_9 = _T_16258 | _T_9530; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16271 = bht_wr_en0[1] & _T_11918; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16275 = _T_16271 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_10 = _T_16275 | _T_9539; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16288 = bht_wr_en0[1] & _T_11935; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16292 = _T_16288 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_11 = _T_16292 | _T_9548; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16305 = bht_wr_en0[1] & _T_11952; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16309 = _T_16305 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_12 = _T_16309 | _T_9557; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16322 = bht_wr_en0[1] & _T_11969; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16326 = _T_16322 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_13 = _T_16326 | _T_9566; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16339 = bht_wr_en0[1] & _T_11986; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16343 = _T_16339 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_14 = _T_16343 | _T_9575; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16356 = bht_wr_en0[1] & _T_12003; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_16360 = _T_16356 & _T_6788; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_15 = _T_16360 | _T_9584; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16377 = _T_16101 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_0 = _T_16377 | _T_9593; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16394 = _T_16118 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_1 = _T_16394 | _T_9602; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16411 = _T_16135 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_2 = _T_16411 | _T_9611; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16428 = _T_16152 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_3 = _T_16428 | _T_9620; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16445 = _T_16169 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_4 = _T_16445 | _T_9629; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16462 = _T_16186 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_5 = _T_16462 | _T_9638; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16479 = _T_16203 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_6 = _T_16479 | _T_9647; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16496 = _T_16220 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_7 = _T_16496 | _T_9656; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16513 = _T_16237 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_8 = _T_16513 | _T_9665; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16530 = _T_16254 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_9 = _T_16530 | _T_9674; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16547 = _T_16271 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_10 = _T_16547 | _T_9683; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16564 = _T_16288 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_11 = _T_16564 | _T_9692; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16581 = _T_16305 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_12 = _T_16581 | _T_9701; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16598 = _T_16322 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_13 = _T_16598 | _T_9710; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16615 = _T_16339 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_14 = _T_16615 | _T_9719; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16632 = _T_16356 & _T_6799; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_15 = _T_16632 | _T_9728; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16649 = _T_16101 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_0 = _T_16649 | _T_9737; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16666 = _T_16118 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_1 = _T_16666 | _T_9746; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16683 = _T_16135 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_2 = _T_16683 | _T_9755; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16700 = _T_16152 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_3 = _T_16700 | _T_9764; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16717 = _T_16169 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_4 = _T_16717 | _T_9773; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16734 = _T_16186 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_5 = _T_16734 | _T_9782; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16751 = _T_16203 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_6 = _T_16751 | _T_9791; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16768 = _T_16220 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_7 = _T_16768 | _T_9800; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16785 = _T_16237 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_8 = _T_16785 | _T_9809; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16802 = _T_16254 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_9 = _T_16802 | _T_9818; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16819 = _T_16271 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_10 = _T_16819 | _T_9827; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16836 = _T_16288 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_11 = _T_16836 | _T_9836; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16853 = _T_16305 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_12 = _T_16853 | _T_9845; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16870 = _T_16322 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_13 = _T_16870 | _T_9854; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16887 = _T_16339 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_14 = _T_16887 | _T_9863; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16904 = _T_16356 & _T_6810; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_15 = _T_16904 | _T_9872; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16921 = _T_16101 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_0 = _T_16921 | _T_9881; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16938 = _T_16118 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_1 = _T_16938 | _T_9890; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16955 = _T_16135 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_2 = _T_16955 | _T_9899; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16972 = _T_16152 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_3 = _T_16972 | _T_9908; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16989 = _T_16169 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_4 = _T_16989 | _T_9917; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17006 = _T_16186 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_5 = _T_17006 | _T_9926; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17023 = _T_16203 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_6 = _T_17023 | _T_9935; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17040 = _T_16220 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_7 = _T_17040 | _T_9944; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17057 = _T_16237 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_8 = _T_17057 | _T_9953; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17074 = _T_16254 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_9 = _T_17074 | _T_9962; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17091 = _T_16271 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_10 = _T_17091 | _T_9971; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17108 = _T_16288 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_11 = _T_17108 | _T_9980; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17125 = _T_16305 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_12 = _T_17125 | _T_9989; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17142 = _T_16322 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_13 = _T_17142 | _T_9998; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17159 = _T_16339 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_14 = _T_17159 | _T_10007; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17176 = _T_16356 & _T_6821; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_15 = _T_17176 | _T_10016; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17193 = _T_16101 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_0 = _T_17193 | _T_10025; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17210 = _T_16118 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_1 = _T_17210 | _T_10034; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17227 = _T_16135 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_2 = _T_17227 | _T_10043; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17244 = _T_16152 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_3 = _T_17244 | _T_10052; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17261 = _T_16169 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_4 = _T_17261 | _T_10061; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17278 = _T_16186 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_5 = _T_17278 | _T_10070; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17295 = _T_16203 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_6 = _T_17295 | _T_10079; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17312 = _T_16220 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_7 = _T_17312 | _T_10088; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17329 = _T_16237 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_8 = _T_17329 | _T_10097; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17346 = _T_16254 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_9 = _T_17346 | _T_10106; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17363 = _T_16271 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_10 = _T_17363 | _T_10115; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17380 = _T_16288 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_11 = _T_17380 | _T_10124; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17397 = _T_16305 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_12 = _T_17397 | _T_10133; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17414 = _T_16322 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_13 = _T_17414 | _T_10142; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17431 = _T_16339 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_14 = _T_17431 | _T_10151; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17448 = _T_16356 & _T_6832; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_15 = _T_17448 | _T_10160; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17465 = _T_16101 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_0 = _T_17465 | _T_10169; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17482 = _T_16118 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_1 = _T_17482 | _T_10178; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17499 = _T_16135 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_2 = _T_17499 | _T_10187; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17516 = _T_16152 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_3 = _T_17516 | _T_10196; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17533 = _T_16169 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_4 = _T_17533 | _T_10205; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17550 = _T_16186 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_5 = _T_17550 | _T_10214; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17567 = _T_16203 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_6 = _T_17567 | _T_10223; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17584 = _T_16220 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_7 = _T_17584 | _T_10232; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17601 = _T_16237 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_8 = _T_17601 | _T_10241; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17618 = _T_16254 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_9 = _T_17618 | _T_10250; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17635 = _T_16271 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_10 = _T_17635 | _T_10259; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17652 = _T_16288 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_11 = _T_17652 | _T_10268; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17669 = _T_16305 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_12 = _T_17669 | _T_10277; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17686 = _T_16322 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_13 = _T_17686 | _T_10286; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17703 = _T_16339 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_14 = _T_17703 | _T_10295; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17720 = _T_16356 & _T_6843; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_15 = _T_17720 | _T_10304; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17737 = _T_16101 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_0 = _T_17737 | _T_10313; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17754 = _T_16118 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_1 = _T_17754 | _T_10322; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17771 = _T_16135 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_2 = _T_17771 | _T_10331; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17788 = _T_16152 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_3 = _T_17788 | _T_10340; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17805 = _T_16169 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_4 = _T_17805 | _T_10349; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17822 = _T_16186 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_5 = _T_17822 | _T_10358; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17839 = _T_16203 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_6 = _T_17839 | _T_10367; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17856 = _T_16220 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_7 = _T_17856 | _T_10376; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17873 = _T_16237 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_8 = _T_17873 | _T_10385; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17890 = _T_16254 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_9 = _T_17890 | _T_10394; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17907 = _T_16271 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_10 = _T_17907 | _T_10403; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17924 = _T_16288 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_11 = _T_17924 | _T_10412; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17941 = _T_16305 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_12 = _T_17941 | _T_10421; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17958 = _T_16322 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_13 = _T_17958 | _T_10430; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17975 = _T_16339 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_14 = _T_17975 | _T_10439; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17992 = _T_16356 & _T_6854; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_15 = _T_17992 | _T_10448; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18009 = _T_16101 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_0 = _T_18009 | _T_10457; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18026 = _T_16118 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_1 = _T_18026 | _T_10466; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18043 = _T_16135 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_2 = _T_18043 | _T_10475; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18060 = _T_16152 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_3 = _T_18060 | _T_10484; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18077 = _T_16169 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_4 = _T_18077 | _T_10493; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18094 = _T_16186 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_5 = _T_18094 | _T_10502; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18111 = _T_16203 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_6 = _T_18111 | _T_10511; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18128 = _T_16220 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_7 = _T_18128 | _T_10520; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18145 = _T_16237 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_8 = _T_18145 | _T_10529; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18162 = _T_16254 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_9 = _T_18162 | _T_10538; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18179 = _T_16271 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_10 = _T_18179 | _T_10547; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18196 = _T_16288 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_11 = _T_18196 | _T_10556; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18213 = _T_16305 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_12 = _T_18213 | _T_10565; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18230 = _T_16322 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_13 = _T_18230 | _T_10574; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18247 = _T_16339 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_14 = _T_18247 | _T_10583; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18264 = _T_16356 & _T_6865; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_15 = _T_18264 | _T_10592; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18281 = _T_16101 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_0 = _T_18281 | _T_10601; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18298 = _T_16118 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_1 = _T_18298 | _T_10610; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18315 = _T_16135 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_2 = _T_18315 | _T_10619; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18332 = _T_16152 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_3 = _T_18332 | _T_10628; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18349 = _T_16169 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_4 = _T_18349 | _T_10637; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18366 = _T_16186 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_5 = _T_18366 | _T_10646; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18383 = _T_16203 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_6 = _T_18383 | _T_10655; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18400 = _T_16220 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_7 = _T_18400 | _T_10664; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18417 = _T_16237 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_8 = _T_18417 | _T_10673; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18434 = _T_16254 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_9 = _T_18434 | _T_10682; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18451 = _T_16271 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_10 = _T_18451 | _T_10691; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18468 = _T_16288 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_11 = _T_18468 | _T_10700; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18485 = _T_16305 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_12 = _T_18485 | _T_10709; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18502 = _T_16322 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_13 = _T_18502 | _T_10718; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18519 = _T_16339 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_14 = _T_18519 | _T_10727; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18536 = _T_16356 & _T_6876; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_15 = _T_18536 | _T_10736; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18553 = _T_16101 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_0 = _T_18553 | _T_10745; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18570 = _T_16118 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_1 = _T_18570 | _T_10754; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18587 = _T_16135 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_2 = _T_18587 | _T_10763; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18604 = _T_16152 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_3 = _T_18604 | _T_10772; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18621 = _T_16169 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_4 = _T_18621 | _T_10781; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18638 = _T_16186 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_5 = _T_18638 | _T_10790; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18655 = _T_16203 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_6 = _T_18655 | _T_10799; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18672 = _T_16220 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_7 = _T_18672 | _T_10808; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18689 = _T_16237 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_8 = _T_18689 | _T_10817; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18706 = _T_16254 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_9 = _T_18706 | _T_10826; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18723 = _T_16271 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_10 = _T_18723 | _T_10835; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18740 = _T_16288 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_11 = _T_18740 | _T_10844; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18757 = _T_16305 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_12 = _T_18757 | _T_10853; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18774 = _T_16322 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_13 = _T_18774 | _T_10862; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18791 = _T_16339 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_14 = _T_18791 | _T_10871; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18808 = _T_16356 & _T_6887; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_15 = _T_18808 | _T_10880; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18825 = _T_16101 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_0 = _T_18825 | _T_10889; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18842 = _T_16118 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_1 = _T_18842 | _T_10898; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18859 = _T_16135 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_2 = _T_18859 | _T_10907; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18876 = _T_16152 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_3 = _T_18876 | _T_10916; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18893 = _T_16169 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_4 = _T_18893 | _T_10925; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18910 = _T_16186 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_5 = _T_18910 | _T_10934; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18927 = _T_16203 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_6 = _T_18927 | _T_10943; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18944 = _T_16220 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_7 = _T_18944 | _T_10952; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18961 = _T_16237 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_8 = _T_18961 | _T_10961; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18978 = _T_16254 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_9 = _T_18978 | _T_10970; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18995 = _T_16271 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_10 = _T_18995 | _T_10979; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19012 = _T_16288 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_11 = _T_19012 | _T_10988; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19029 = _T_16305 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_12 = _T_19029 | _T_10997; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19046 = _T_16322 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_13 = _T_19046 | _T_11006; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19063 = _T_16339 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_14 = _T_19063 | _T_11015; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19080 = _T_16356 & _T_6898; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_15 = _T_19080 | _T_11024; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19097 = _T_16101 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_0 = _T_19097 | _T_11033; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19114 = _T_16118 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_1 = _T_19114 | _T_11042; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19131 = _T_16135 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_2 = _T_19131 | _T_11051; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19148 = _T_16152 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_3 = _T_19148 | _T_11060; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19165 = _T_16169 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_4 = _T_19165 | _T_11069; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19182 = _T_16186 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_5 = _T_19182 | _T_11078; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19199 = _T_16203 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_6 = _T_19199 | _T_11087; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19216 = _T_16220 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_7 = _T_19216 | _T_11096; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19233 = _T_16237 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_8 = _T_19233 | _T_11105; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19250 = _T_16254 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_9 = _T_19250 | _T_11114; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19267 = _T_16271 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_10 = _T_19267 | _T_11123; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19284 = _T_16288 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_11 = _T_19284 | _T_11132; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19301 = _T_16305 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_12 = _T_19301 | _T_11141; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19318 = _T_16322 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_13 = _T_19318 | _T_11150; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19335 = _T_16339 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_14 = _T_19335 | _T_11159; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19352 = _T_16356 & _T_6909; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_15 = _T_19352 | _T_11168; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19369 = _T_16101 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_0 = _T_19369 | _T_11177; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19386 = _T_16118 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_1 = _T_19386 | _T_11186; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19403 = _T_16135 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_2 = _T_19403 | _T_11195; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19420 = _T_16152 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_3 = _T_19420 | _T_11204; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19437 = _T_16169 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_4 = _T_19437 | _T_11213; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19454 = _T_16186 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_5 = _T_19454 | _T_11222; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19471 = _T_16203 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_6 = _T_19471 | _T_11231; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19488 = _T_16220 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_7 = _T_19488 | _T_11240; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19505 = _T_16237 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_8 = _T_19505 | _T_11249; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19522 = _T_16254 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_9 = _T_19522 | _T_11258; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19539 = _T_16271 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_10 = _T_19539 | _T_11267; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19556 = _T_16288 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_11 = _T_19556 | _T_11276; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19573 = _T_16305 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_12 = _T_19573 | _T_11285; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19590 = _T_16322 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_13 = _T_19590 | _T_11294; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19607 = _T_16339 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_14 = _T_19607 | _T_11303; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19624 = _T_16356 & _T_6920; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_15 = _T_19624 | _T_11312; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19641 = _T_16101 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_0 = _T_19641 | _T_11321; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19658 = _T_16118 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_1 = _T_19658 | _T_11330; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19675 = _T_16135 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_2 = _T_19675 | _T_11339; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19692 = _T_16152 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_3 = _T_19692 | _T_11348; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19709 = _T_16169 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_4 = _T_19709 | _T_11357; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19726 = _T_16186 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_5 = _T_19726 | _T_11366; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19743 = _T_16203 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_6 = _T_19743 | _T_11375; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19760 = _T_16220 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_7 = _T_19760 | _T_11384; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19777 = _T_16237 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_8 = _T_19777 | _T_11393; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19794 = _T_16254 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_9 = _T_19794 | _T_11402; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19811 = _T_16271 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_10 = _T_19811 | _T_11411; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19828 = _T_16288 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_11 = _T_19828 | _T_11420; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19845 = _T_16305 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_12 = _T_19845 | _T_11429; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19862 = _T_16322 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_13 = _T_19862 | _T_11438; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19879 = _T_16339 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_14 = _T_19879 | _T_11447; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19896 = _T_16356 & _T_6931; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_15 = _T_19896 | _T_11456; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19913 = _T_16101 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_0 = _T_19913 | _T_11465; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19930 = _T_16118 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_1 = _T_19930 | _T_11474; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19947 = _T_16135 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_2 = _T_19947 | _T_11483; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19964 = _T_16152 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_3 = _T_19964 | _T_11492; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19981 = _T_16169 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_4 = _T_19981 | _T_11501; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19998 = _T_16186 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_5 = _T_19998 | _T_11510; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20015 = _T_16203 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_6 = _T_20015 | _T_11519; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20032 = _T_16220 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_7 = _T_20032 | _T_11528; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20049 = _T_16237 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_8 = _T_20049 | _T_11537; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20066 = _T_16254 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_9 = _T_20066 | _T_11546; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20083 = _T_16271 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_10 = _T_20083 | _T_11555; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20100 = _T_16288 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_11 = _T_20100 | _T_11564; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20117 = _T_16305 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_12 = _T_20117 | _T_11573; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20134 = _T_16322 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_13 = _T_20134 | _T_11582; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20151 = _T_16339 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_14 = _T_20151 | _T_11591; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20168 = _T_16356 & _T_6942; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_15 = _T_20168 | _T_11600; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20185 = _T_16101 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_0 = _T_20185 | _T_11609; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20202 = _T_16118 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_1 = _T_20202 | _T_11618; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20219 = _T_16135 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_2 = _T_20219 | _T_11627; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20236 = _T_16152 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_3 = _T_20236 | _T_11636; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20253 = _T_16169 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_4 = _T_20253 | _T_11645; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20270 = _T_16186 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_5 = _T_20270 | _T_11654; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20287 = _T_16203 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_6 = _T_20287 | _T_11663; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20304 = _T_16220 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_7 = _T_20304 | _T_11672; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20321 = _T_16237 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_8 = _T_20321 | _T_11681; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20338 = _T_16254 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_9 = _T_20338 | _T_11690; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20355 = _T_16271 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_10 = _T_20355 | _T_11699; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20372 = _T_16288 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_11 = _T_20372 | _T_11708; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20389 = _T_16305 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_12 = _T_20389 | _T_11717; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20406 = _T_16322 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_13 = _T_20406 | _T_11726; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20423 = _T_16339 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_14 = _T_20423 | _T_11735; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_20440 = _T_16356 & _T_6953; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_15 = _T_20440 | _T_11744; // @[ifu_bp_ctl.scala 526:223]
  rvclkhdr rvclkhdr ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en)
  );
  rvclkhdr rvclkhdr_20 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en)
  );
  rvclkhdr rvclkhdr_21 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en)
  );
  rvclkhdr rvclkhdr_22 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en)
  );
  rvclkhdr rvclkhdr_23 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en)
  );
  rvclkhdr rvclkhdr_24 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en)
  );
  rvclkhdr rvclkhdr_25 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en)
  );
  rvclkhdr rvclkhdr_26 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en)
  );
  rvclkhdr rvclkhdr_27 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en)
  );
  rvclkhdr rvclkhdr_28 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en)
  );
  rvclkhdr rvclkhdr_29 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en)
  );
  rvclkhdr rvclkhdr_30 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en)
  );
  rvclkhdr rvclkhdr_31 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en)
  );
  rvclkhdr rvclkhdr_32 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en)
  );
  rvclkhdr rvclkhdr_33 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en)
  );
  rvclkhdr rvclkhdr_34 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en)
  );
  rvclkhdr rvclkhdr_35 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en)
  );
  rvclkhdr rvclkhdr_36 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en)
  );
  rvclkhdr rvclkhdr_37 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en)
  );
  rvclkhdr rvclkhdr_38 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en)
  );
  rvclkhdr rvclkhdr_39 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en)
  );
  rvclkhdr rvclkhdr_40 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en)
  );
  rvclkhdr rvclkhdr_41 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en)
  );
  rvclkhdr rvclkhdr_42 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en)
  );
  rvclkhdr rvclkhdr_43 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en)
  );
  rvclkhdr rvclkhdr_44 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en)
  );
  rvclkhdr rvclkhdr_45 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en)
  );
  rvclkhdr rvclkhdr_46 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en)
  );
  rvclkhdr rvclkhdr_47 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en)
  );
  rvclkhdr rvclkhdr_48 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en)
  );
  rvclkhdr rvclkhdr_49 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en)
  );
  rvclkhdr rvclkhdr_50 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en)
  );
  rvclkhdr rvclkhdr_51 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en)
  );
  rvclkhdr rvclkhdr_52 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en)
  );
  rvclkhdr rvclkhdr_53 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en)
  );
  rvclkhdr rvclkhdr_54 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en)
  );
  rvclkhdr rvclkhdr_55 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en)
  );
  rvclkhdr rvclkhdr_56 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en)
  );
  rvclkhdr rvclkhdr_57 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en)
  );
  rvclkhdr rvclkhdr_58 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en)
  );
  rvclkhdr rvclkhdr_59 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en)
  );
  rvclkhdr rvclkhdr_60 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en)
  );
  rvclkhdr rvclkhdr_61 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en)
  );
  rvclkhdr rvclkhdr_62 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en)
  );
  rvclkhdr rvclkhdr_63 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en)
  );
  rvclkhdr rvclkhdr_64 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en)
  );
  rvclkhdr rvclkhdr_65 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en)
  );
  rvclkhdr rvclkhdr_66 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en)
  );
  rvclkhdr rvclkhdr_67 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en)
  );
  rvclkhdr rvclkhdr_68 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en)
  );
  rvclkhdr rvclkhdr_69 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en)
  );
  rvclkhdr rvclkhdr_70 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en)
  );
  rvclkhdr rvclkhdr_71 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en)
  );
  rvclkhdr rvclkhdr_72 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en)
  );
  rvclkhdr rvclkhdr_73 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en)
  );
  rvclkhdr rvclkhdr_74 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en)
  );
  rvclkhdr rvclkhdr_75 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en)
  );
  rvclkhdr rvclkhdr_76 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en)
  );
  rvclkhdr rvclkhdr_77 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en)
  );
  rvclkhdr rvclkhdr_78 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en)
  );
  rvclkhdr rvclkhdr_79 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en)
  );
  rvclkhdr rvclkhdr_80 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en)
  );
  rvclkhdr rvclkhdr_81 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en)
  );
  rvclkhdr rvclkhdr_82 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en)
  );
  rvclkhdr rvclkhdr_83 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en)
  );
  rvclkhdr rvclkhdr_84 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en)
  );
  rvclkhdr rvclkhdr_85 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en)
  );
  rvclkhdr rvclkhdr_86 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en)
  );
  rvclkhdr rvclkhdr_87 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en)
  );
  rvclkhdr rvclkhdr_88 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en)
  );
  rvclkhdr rvclkhdr_89 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en)
  );
  rvclkhdr rvclkhdr_90 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en)
  );
  rvclkhdr rvclkhdr_91 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en)
  );
  rvclkhdr rvclkhdr_92 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en)
  );
  rvclkhdr rvclkhdr_93 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en)
  );
  rvclkhdr rvclkhdr_94 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_94_io_clk),
    .io_en(rvclkhdr_94_io_en)
  );
  rvclkhdr rvclkhdr_95 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_95_io_clk),
    .io_en(rvclkhdr_95_io_en)
  );
  rvclkhdr rvclkhdr_96 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_96_io_clk),
    .io_en(rvclkhdr_96_io_en)
  );
  rvclkhdr rvclkhdr_97 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_97_io_clk),
    .io_en(rvclkhdr_97_io_en)
  );
  rvclkhdr rvclkhdr_98 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_98_io_clk),
    .io_en(rvclkhdr_98_io_en)
  );
  rvclkhdr rvclkhdr_99 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_99_io_clk),
    .io_en(rvclkhdr_99_io_en)
  );
  rvclkhdr rvclkhdr_100 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_100_io_clk),
    .io_en(rvclkhdr_100_io_en)
  );
  rvclkhdr rvclkhdr_101 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_101_io_clk),
    .io_en(rvclkhdr_101_io_en)
  );
  rvclkhdr rvclkhdr_102 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_102_io_clk),
    .io_en(rvclkhdr_102_io_en)
  );
  rvclkhdr rvclkhdr_103 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_103_io_clk),
    .io_en(rvclkhdr_103_io_en)
  );
  rvclkhdr rvclkhdr_104 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_104_io_clk),
    .io_en(rvclkhdr_104_io_en)
  );
  rvclkhdr rvclkhdr_105 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_105_io_clk),
    .io_en(rvclkhdr_105_io_en)
  );
  rvclkhdr rvclkhdr_106 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_106_io_clk),
    .io_en(rvclkhdr_106_io_en)
  );
  rvclkhdr rvclkhdr_107 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_107_io_clk),
    .io_en(rvclkhdr_107_io_en)
  );
  rvclkhdr rvclkhdr_108 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_108_io_clk),
    .io_en(rvclkhdr_108_io_en)
  );
  rvclkhdr rvclkhdr_109 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_109_io_clk),
    .io_en(rvclkhdr_109_io_en)
  );
  rvclkhdr rvclkhdr_110 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_110_io_clk),
    .io_en(rvclkhdr_110_io_en)
  );
  rvclkhdr rvclkhdr_111 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_111_io_clk),
    .io_en(rvclkhdr_111_io_en)
  );
  rvclkhdr rvclkhdr_112 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_112_io_clk),
    .io_en(rvclkhdr_112_io_en)
  );
  rvclkhdr rvclkhdr_113 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_113_io_clk),
    .io_en(rvclkhdr_113_io_en)
  );
  rvclkhdr rvclkhdr_114 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_114_io_clk),
    .io_en(rvclkhdr_114_io_en)
  );
  rvclkhdr rvclkhdr_115 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_115_io_clk),
    .io_en(rvclkhdr_115_io_en)
  );
  rvclkhdr rvclkhdr_116 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_116_io_clk),
    .io_en(rvclkhdr_116_io_en)
  );
  rvclkhdr rvclkhdr_117 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_117_io_clk),
    .io_en(rvclkhdr_117_io_en)
  );
  rvclkhdr rvclkhdr_118 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_118_io_clk),
    .io_en(rvclkhdr_118_io_en)
  );
  rvclkhdr rvclkhdr_119 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_119_io_clk),
    .io_en(rvclkhdr_119_io_en)
  );
  rvclkhdr rvclkhdr_120 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_120_io_clk),
    .io_en(rvclkhdr_120_io_en)
  );
  rvclkhdr rvclkhdr_121 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_121_io_clk),
    .io_en(rvclkhdr_121_io_en)
  );
  rvclkhdr rvclkhdr_122 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_122_io_clk),
    .io_en(rvclkhdr_122_io_en)
  );
  rvclkhdr rvclkhdr_123 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_123_io_clk),
    .io_en(rvclkhdr_123_io_en)
  );
  rvclkhdr rvclkhdr_124 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_124_io_clk),
    .io_en(rvclkhdr_124_io_en)
  );
  rvclkhdr rvclkhdr_125 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_125_io_clk),
    .io_en(rvclkhdr_125_io_en)
  );
  rvclkhdr rvclkhdr_126 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_126_io_clk),
    .io_en(rvclkhdr_126_io_en)
  );
  rvclkhdr rvclkhdr_127 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_127_io_clk),
    .io_en(rvclkhdr_127_io_en)
  );
  rvclkhdr rvclkhdr_128 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_128_io_clk),
    .io_en(rvclkhdr_128_io_en)
  );
  rvclkhdr rvclkhdr_129 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_129_io_clk),
    .io_en(rvclkhdr_129_io_en)
  );
  rvclkhdr rvclkhdr_130 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_130_io_clk),
    .io_en(rvclkhdr_130_io_en)
  );
  rvclkhdr rvclkhdr_131 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_131_io_clk),
    .io_en(rvclkhdr_131_io_en)
  );
  rvclkhdr rvclkhdr_132 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_132_io_clk),
    .io_en(rvclkhdr_132_io_en)
  );
  rvclkhdr rvclkhdr_133 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_133_io_clk),
    .io_en(rvclkhdr_133_io_en)
  );
  rvclkhdr rvclkhdr_134 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_134_io_clk),
    .io_en(rvclkhdr_134_io_en)
  );
  rvclkhdr rvclkhdr_135 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_135_io_clk),
    .io_en(rvclkhdr_135_io_en)
  );
  rvclkhdr rvclkhdr_136 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_136_io_clk),
    .io_en(rvclkhdr_136_io_en)
  );
  rvclkhdr rvclkhdr_137 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_137_io_clk),
    .io_en(rvclkhdr_137_io_en)
  );
  rvclkhdr rvclkhdr_138 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_138_io_clk),
    .io_en(rvclkhdr_138_io_en)
  );
  rvclkhdr rvclkhdr_139 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_139_io_clk),
    .io_en(rvclkhdr_139_io_en)
  );
  rvclkhdr rvclkhdr_140 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_140_io_clk),
    .io_en(rvclkhdr_140_io_en)
  );
  rvclkhdr rvclkhdr_141 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_141_io_clk),
    .io_en(rvclkhdr_141_io_en)
  );
  rvclkhdr rvclkhdr_142 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_142_io_clk),
    .io_en(rvclkhdr_142_io_en)
  );
  rvclkhdr rvclkhdr_143 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_143_io_clk),
    .io_en(rvclkhdr_143_io_en)
  );
  rvclkhdr rvclkhdr_144 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_144_io_clk),
    .io_en(rvclkhdr_144_io_en)
  );
  rvclkhdr rvclkhdr_145 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_145_io_clk),
    .io_en(rvclkhdr_145_io_en)
  );
  rvclkhdr rvclkhdr_146 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_146_io_clk),
    .io_en(rvclkhdr_146_io_en)
  );
  rvclkhdr rvclkhdr_147 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_147_io_clk),
    .io_en(rvclkhdr_147_io_en)
  );
  rvclkhdr rvclkhdr_148 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_148_io_clk),
    .io_en(rvclkhdr_148_io_en)
  );
  rvclkhdr rvclkhdr_149 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_149_io_clk),
    .io_en(rvclkhdr_149_io_en)
  );
  rvclkhdr rvclkhdr_150 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_150_io_clk),
    .io_en(rvclkhdr_150_io_en)
  );
  rvclkhdr rvclkhdr_151 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_151_io_clk),
    .io_en(rvclkhdr_151_io_en)
  );
  rvclkhdr rvclkhdr_152 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_152_io_clk),
    .io_en(rvclkhdr_152_io_en)
  );
  rvclkhdr rvclkhdr_153 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_153_io_clk),
    .io_en(rvclkhdr_153_io_en)
  );
  rvclkhdr rvclkhdr_154 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_154_io_clk),
    .io_en(rvclkhdr_154_io_en)
  );
  rvclkhdr rvclkhdr_155 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_155_io_clk),
    .io_en(rvclkhdr_155_io_en)
  );
  rvclkhdr rvclkhdr_156 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_156_io_clk),
    .io_en(rvclkhdr_156_io_en)
  );
  rvclkhdr rvclkhdr_157 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_157_io_clk),
    .io_en(rvclkhdr_157_io_en)
  );
  rvclkhdr rvclkhdr_158 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_158_io_clk),
    .io_en(rvclkhdr_158_io_en)
  );
  rvclkhdr rvclkhdr_159 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_159_io_clk),
    .io_en(rvclkhdr_159_io_en)
  );
  rvclkhdr rvclkhdr_160 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_160_io_clk),
    .io_en(rvclkhdr_160_io_en)
  );
  rvclkhdr rvclkhdr_161 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_161_io_clk),
    .io_en(rvclkhdr_161_io_en)
  );
  rvclkhdr rvclkhdr_162 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_162_io_clk),
    .io_en(rvclkhdr_162_io_en)
  );
  rvclkhdr rvclkhdr_163 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_163_io_clk),
    .io_en(rvclkhdr_163_io_en)
  );
  rvclkhdr rvclkhdr_164 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_164_io_clk),
    .io_en(rvclkhdr_164_io_en)
  );
  rvclkhdr rvclkhdr_165 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_165_io_clk),
    .io_en(rvclkhdr_165_io_en)
  );
  rvclkhdr rvclkhdr_166 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_166_io_clk),
    .io_en(rvclkhdr_166_io_en)
  );
  rvclkhdr rvclkhdr_167 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_167_io_clk),
    .io_en(rvclkhdr_167_io_en)
  );
  rvclkhdr rvclkhdr_168 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_168_io_clk),
    .io_en(rvclkhdr_168_io_en)
  );
  rvclkhdr rvclkhdr_169 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_169_io_clk),
    .io_en(rvclkhdr_169_io_en)
  );
  rvclkhdr rvclkhdr_170 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_170_io_clk),
    .io_en(rvclkhdr_170_io_en)
  );
  rvclkhdr rvclkhdr_171 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_171_io_clk),
    .io_en(rvclkhdr_171_io_en)
  );
  rvclkhdr rvclkhdr_172 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_172_io_clk),
    .io_en(rvclkhdr_172_io_en)
  );
  rvclkhdr rvclkhdr_173 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_173_io_clk),
    .io_en(rvclkhdr_173_io_en)
  );
  rvclkhdr rvclkhdr_174 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_174_io_clk),
    .io_en(rvclkhdr_174_io_en)
  );
  rvclkhdr rvclkhdr_175 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_175_io_clk),
    .io_en(rvclkhdr_175_io_en)
  );
  rvclkhdr rvclkhdr_176 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_176_io_clk),
    .io_en(rvclkhdr_176_io_en)
  );
  rvclkhdr rvclkhdr_177 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_177_io_clk),
    .io_en(rvclkhdr_177_io_en)
  );
  rvclkhdr rvclkhdr_178 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_178_io_clk),
    .io_en(rvclkhdr_178_io_en)
  );
  rvclkhdr rvclkhdr_179 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_179_io_clk),
    .io_en(rvclkhdr_179_io_en)
  );
  rvclkhdr rvclkhdr_180 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_180_io_clk),
    .io_en(rvclkhdr_180_io_en)
  );
  rvclkhdr rvclkhdr_181 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_181_io_clk),
    .io_en(rvclkhdr_181_io_en)
  );
  rvclkhdr rvclkhdr_182 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_182_io_clk),
    .io_en(rvclkhdr_182_io_en)
  );
  rvclkhdr rvclkhdr_183 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_183_io_clk),
    .io_en(rvclkhdr_183_io_en)
  );
  rvclkhdr rvclkhdr_184 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_184_io_clk),
    .io_en(rvclkhdr_184_io_en)
  );
  rvclkhdr rvclkhdr_185 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_185_io_clk),
    .io_en(rvclkhdr_185_io_en)
  );
  rvclkhdr rvclkhdr_186 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_186_io_clk),
    .io_en(rvclkhdr_186_io_en)
  );
  rvclkhdr rvclkhdr_187 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_187_io_clk),
    .io_en(rvclkhdr_187_io_en)
  );
  rvclkhdr rvclkhdr_188 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_188_io_clk),
    .io_en(rvclkhdr_188_io_en)
  );
  rvclkhdr rvclkhdr_189 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_189_io_clk),
    .io_en(rvclkhdr_189_io_en)
  );
  rvclkhdr rvclkhdr_190 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_190_io_clk),
    .io_en(rvclkhdr_190_io_en)
  );
  rvclkhdr rvclkhdr_191 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_191_io_clk),
    .io_en(rvclkhdr_191_io_en)
  );
  rvclkhdr rvclkhdr_192 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_192_io_clk),
    .io_en(rvclkhdr_192_io_en)
  );
  rvclkhdr rvclkhdr_193 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_193_io_clk),
    .io_en(rvclkhdr_193_io_en)
  );
  rvclkhdr rvclkhdr_194 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_194_io_clk),
    .io_en(rvclkhdr_194_io_en)
  );
  rvclkhdr rvclkhdr_195 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_195_io_clk),
    .io_en(rvclkhdr_195_io_en)
  );
  rvclkhdr rvclkhdr_196 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_196_io_clk),
    .io_en(rvclkhdr_196_io_en)
  );
  rvclkhdr rvclkhdr_197 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_197_io_clk),
    .io_en(rvclkhdr_197_io_en)
  );
  rvclkhdr rvclkhdr_198 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_198_io_clk),
    .io_en(rvclkhdr_198_io_en)
  );
  rvclkhdr rvclkhdr_199 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_199_io_clk),
    .io_en(rvclkhdr_199_io_en)
  );
  rvclkhdr rvclkhdr_200 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_200_io_clk),
    .io_en(rvclkhdr_200_io_en)
  );
  rvclkhdr rvclkhdr_201 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_201_io_clk),
    .io_en(rvclkhdr_201_io_en)
  );
  rvclkhdr rvclkhdr_202 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_202_io_clk),
    .io_en(rvclkhdr_202_io_en)
  );
  rvclkhdr rvclkhdr_203 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_203_io_clk),
    .io_en(rvclkhdr_203_io_en)
  );
  rvclkhdr rvclkhdr_204 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_204_io_clk),
    .io_en(rvclkhdr_204_io_en)
  );
  rvclkhdr rvclkhdr_205 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_205_io_clk),
    .io_en(rvclkhdr_205_io_en)
  );
  rvclkhdr rvclkhdr_206 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_206_io_clk),
    .io_en(rvclkhdr_206_io_en)
  );
  rvclkhdr rvclkhdr_207 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_207_io_clk),
    .io_en(rvclkhdr_207_io_en)
  );
  rvclkhdr rvclkhdr_208 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_208_io_clk),
    .io_en(rvclkhdr_208_io_en)
  );
  rvclkhdr rvclkhdr_209 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_209_io_clk),
    .io_en(rvclkhdr_209_io_en)
  );
  rvclkhdr rvclkhdr_210 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_210_io_clk),
    .io_en(rvclkhdr_210_io_en)
  );
  rvclkhdr rvclkhdr_211 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_211_io_clk),
    .io_en(rvclkhdr_211_io_en)
  );
  rvclkhdr rvclkhdr_212 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_212_io_clk),
    .io_en(rvclkhdr_212_io_en)
  );
  rvclkhdr rvclkhdr_213 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_213_io_clk),
    .io_en(rvclkhdr_213_io_en)
  );
  rvclkhdr rvclkhdr_214 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_214_io_clk),
    .io_en(rvclkhdr_214_io_en)
  );
  rvclkhdr rvclkhdr_215 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_215_io_clk),
    .io_en(rvclkhdr_215_io_en)
  );
  rvclkhdr rvclkhdr_216 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_216_io_clk),
    .io_en(rvclkhdr_216_io_en)
  );
  rvclkhdr rvclkhdr_217 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_217_io_clk),
    .io_en(rvclkhdr_217_io_en)
  );
  rvclkhdr rvclkhdr_218 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_218_io_clk),
    .io_en(rvclkhdr_218_io_en)
  );
  rvclkhdr rvclkhdr_219 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_219_io_clk),
    .io_en(rvclkhdr_219_io_en)
  );
  rvclkhdr rvclkhdr_220 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_220_io_clk),
    .io_en(rvclkhdr_220_io_en)
  );
  rvclkhdr rvclkhdr_221 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_221_io_clk),
    .io_en(rvclkhdr_221_io_en)
  );
  rvclkhdr rvclkhdr_222 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_222_io_clk),
    .io_en(rvclkhdr_222_io_en)
  );
  rvclkhdr rvclkhdr_223 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_223_io_clk),
    .io_en(rvclkhdr_223_io_en)
  );
  rvclkhdr rvclkhdr_224 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_224_io_clk),
    .io_en(rvclkhdr_224_io_en)
  );
  rvclkhdr rvclkhdr_225 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_225_io_clk),
    .io_en(rvclkhdr_225_io_en)
  );
  rvclkhdr rvclkhdr_226 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_226_io_clk),
    .io_en(rvclkhdr_226_io_en)
  );
  rvclkhdr rvclkhdr_227 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_227_io_clk),
    .io_en(rvclkhdr_227_io_en)
  );
  rvclkhdr rvclkhdr_228 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_228_io_clk),
    .io_en(rvclkhdr_228_io_en)
  );
  rvclkhdr rvclkhdr_229 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_229_io_clk),
    .io_en(rvclkhdr_229_io_en)
  );
  rvclkhdr rvclkhdr_230 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_230_io_clk),
    .io_en(rvclkhdr_230_io_en)
  );
  rvclkhdr rvclkhdr_231 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_231_io_clk),
    .io_en(rvclkhdr_231_io_en)
  );
  rvclkhdr rvclkhdr_232 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_232_io_clk),
    .io_en(rvclkhdr_232_io_en)
  );
  rvclkhdr rvclkhdr_233 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_233_io_clk),
    .io_en(rvclkhdr_233_io_en)
  );
  rvclkhdr rvclkhdr_234 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_234_io_clk),
    .io_en(rvclkhdr_234_io_en)
  );
  rvclkhdr rvclkhdr_235 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_235_io_clk),
    .io_en(rvclkhdr_235_io_en)
  );
  rvclkhdr rvclkhdr_236 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_236_io_clk),
    .io_en(rvclkhdr_236_io_en)
  );
  rvclkhdr rvclkhdr_237 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_237_io_clk),
    .io_en(rvclkhdr_237_io_en)
  );
  rvclkhdr rvclkhdr_238 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_238_io_clk),
    .io_en(rvclkhdr_238_io_en)
  );
  rvclkhdr rvclkhdr_239 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_239_io_clk),
    .io_en(rvclkhdr_239_io_en)
  );
  rvclkhdr rvclkhdr_240 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_240_io_clk),
    .io_en(rvclkhdr_240_io_en)
  );
  rvclkhdr rvclkhdr_241 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_241_io_clk),
    .io_en(rvclkhdr_241_io_en)
  );
  rvclkhdr rvclkhdr_242 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_242_io_clk),
    .io_en(rvclkhdr_242_io_en)
  );
  rvclkhdr rvclkhdr_243 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_243_io_clk),
    .io_en(rvclkhdr_243_io_en)
  );
  rvclkhdr rvclkhdr_244 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_244_io_clk),
    .io_en(rvclkhdr_244_io_en)
  );
  rvclkhdr rvclkhdr_245 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_245_io_clk),
    .io_en(rvclkhdr_245_io_en)
  );
  rvclkhdr rvclkhdr_246 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_246_io_clk),
    .io_en(rvclkhdr_246_io_en)
  );
  rvclkhdr rvclkhdr_247 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_247_io_clk),
    .io_en(rvclkhdr_247_io_en)
  );
  rvclkhdr rvclkhdr_248 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_248_io_clk),
    .io_en(rvclkhdr_248_io_en)
  );
  rvclkhdr rvclkhdr_249 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_249_io_clk),
    .io_en(rvclkhdr_249_io_en)
  );
  rvclkhdr rvclkhdr_250 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_250_io_clk),
    .io_en(rvclkhdr_250_io_en)
  );
  rvclkhdr rvclkhdr_251 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_251_io_clk),
    .io_en(rvclkhdr_251_io_en)
  );
  rvclkhdr rvclkhdr_252 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_252_io_clk),
    .io_en(rvclkhdr_252_io_en)
  );
  rvclkhdr rvclkhdr_253 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_253_io_clk),
    .io_en(rvclkhdr_253_io_en)
  );
  rvclkhdr rvclkhdr_254 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_254_io_clk),
    .io_en(rvclkhdr_254_io_en)
  );
  rvclkhdr rvclkhdr_255 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_255_io_clk),
    .io_en(rvclkhdr_255_io_en)
  );
  rvclkhdr rvclkhdr_256 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_256_io_clk),
    .io_en(rvclkhdr_256_io_en)
  );
  rvclkhdr rvclkhdr_257 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_257_io_clk),
    .io_en(rvclkhdr_257_io_en)
  );
  rvclkhdr rvclkhdr_258 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_258_io_clk),
    .io_en(rvclkhdr_258_io_en)
  );
  rvclkhdr rvclkhdr_259 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_259_io_clk),
    .io_en(rvclkhdr_259_io_en)
  );
  rvclkhdr rvclkhdr_260 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_260_io_clk),
    .io_en(rvclkhdr_260_io_en)
  );
  rvclkhdr rvclkhdr_261 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_261_io_clk),
    .io_en(rvclkhdr_261_io_en)
  );
  rvclkhdr rvclkhdr_262 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_262_io_clk),
    .io_en(rvclkhdr_262_io_en)
  );
  rvclkhdr rvclkhdr_263 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_263_io_clk),
    .io_en(rvclkhdr_263_io_en)
  );
  rvclkhdr rvclkhdr_264 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_264_io_clk),
    .io_en(rvclkhdr_264_io_en)
  );
  rvclkhdr rvclkhdr_265 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_265_io_clk),
    .io_en(rvclkhdr_265_io_en)
  );
  rvclkhdr rvclkhdr_266 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_266_io_clk),
    .io_en(rvclkhdr_266_io_en)
  );
  rvclkhdr rvclkhdr_267 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_267_io_clk),
    .io_en(rvclkhdr_267_io_en)
  );
  rvclkhdr rvclkhdr_268 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_268_io_clk),
    .io_en(rvclkhdr_268_io_en)
  );
  rvclkhdr rvclkhdr_269 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_269_io_clk),
    .io_en(rvclkhdr_269_io_en)
  );
  rvclkhdr rvclkhdr_270 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_270_io_clk),
    .io_en(rvclkhdr_270_io_en)
  );
  rvclkhdr rvclkhdr_271 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_271_io_clk),
    .io_en(rvclkhdr_271_io_en)
  );
  rvclkhdr rvclkhdr_272 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_272_io_clk),
    .io_en(rvclkhdr_272_io_en)
  );
  rvclkhdr rvclkhdr_273 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_273_io_clk),
    .io_en(rvclkhdr_273_io_en)
  );
  rvclkhdr rvclkhdr_274 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_274_io_clk),
    .io_en(rvclkhdr_274_io_en)
  );
  rvclkhdr rvclkhdr_275 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_275_io_clk),
    .io_en(rvclkhdr_275_io_en)
  );
  rvclkhdr rvclkhdr_276 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_276_io_clk),
    .io_en(rvclkhdr_276_io_en)
  );
  rvclkhdr rvclkhdr_277 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_277_io_clk),
    .io_en(rvclkhdr_277_io_en)
  );
  rvclkhdr rvclkhdr_278 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_278_io_clk),
    .io_en(rvclkhdr_278_io_en)
  );
  rvclkhdr rvclkhdr_279 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_279_io_clk),
    .io_en(rvclkhdr_279_io_en)
  );
  rvclkhdr rvclkhdr_280 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_280_io_clk),
    .io_en(rvclkhdr_280_io_en)
  );
  rvclkhdr rvclkhdr_281 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_281_io_clk),
    .io_en(rvclkhdr_281_io_en)
  );
  rvclkhdr rvclkhdr_282 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_282_io_clk),
    .io_en(rvclkhdr_282_io_en)
  );
  rvclkhdr rvclkhdr_283 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_283_io_clk),
    .io_en(rvclkhdr_283_io_en)
  );
  rvclkhdr rvclkhdr_284 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_284_io_clk),
    .io_en(rvclkhdr_284_io_en)
  );
  rvclkhdr rvclkhdr_285 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_285_io_clk),
    .io_en(rvclkhdr_285_io_en)
  );
  rvclkhdr rvclkhdr_286 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_286_io_clk),
    .io_en(rvclkhdr_286_io_en)
  );
  rvclkhdr rvclkhdr_287 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_287_io_clk),
    .io_en(rvclkhdr_287_io_en)
  );
  rvclkhdr rvclkhdr_288 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_288_io_clk),
    .io_en(rvclkhdr_288_io_en)
  );
  rvclkhdr rvclkhdr_289 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_289_io_clk),
    .io_en(rvclkhdr_289_io_en)
  );
  rvclkhdr rvclkhdr_290 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_290_io_clk),
    .io_en(rvclkhdr_290_io_en)
  );
  rvclkhdr rvclkhdr_291 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_291_io_clk),
    .io_en(rvclkhdr_291_io_en)
  );
  rvclkhdr rvclkhdr_292 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_292_io_clk),
    .io_en(rvclkhdr_292_io_en)
  );
  rvclkhdr rvclkhdr_293 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_293_io_clk),
    .io_en(rvclkhdr_293_io_en)
  );
  rvclkhdr rvclkhdr_294 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_294_io_clk),
    .io_en(rvclkhdr_294_io_en)
  );
  rvclkhdr rvclkhdr_295 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_295_io_clk),
    .io_en(rvclkhdr_295_io_en)
  );
  rvclkhdr rvclkhdr_296 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_296_io_clk),
    .io_en(rvclkhdr_296_io_en)
  );
  rvclkhdr rvclkhdr_297 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_297_io_clk),
    .io_en(rvclkhdr_297_io_en)
  );
  rvclkhdr rvclkhdr_298 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_298_io_clk),
    .io_en(rvclkhdr_298_io_en)
  );
  rvclkhdr rvclkhdr_299 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_299_io_clk),
    .io_en(rvclkhdr_299_io_en)
  );
  rvclkhdr rvclkhdr_300 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_300_io_clk),
    .io_en(rvclkhdr_300_io_en)
  );
  rvclkhdr rvclkhdr_301 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_301_io_clk),
    .io_en(rvclkhdr_301_io_en)
  );
  rvclkhdr rvclkhdr_302 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_302_io_clk),
    .io_en(rvclkhdr_302_io_en)
  );
  rvclkhdr rvclkhdr_303 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_303_io_clk),
    .io_en(rvclkhdr_303_io_en)
  );
  rvclkhdr rvclkhdr_304 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_304_io_clk),
    .io_en(rvclkhdr_304_io_en)
  );
  rvclkhdr rvclkhdr_305 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_305_io_clk),
    .io_en(rvclkhdr_305_io_en)
  );
  rvclkhdr rvclkhdr_306 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_306_io_clk),
    .io_en(rvclkhdr_306_io_en)
  );
  rvclkhdr rvclkhdr_307 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_307_io_clk),
    .io_en(rvclkhdr_307_io_en)
  );
  rvclkhdr rvclkhdr_308 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_308_io_clk),
    .io_en(rvclkhdr_308_io_en)
  );
  rvclkhdr rvclkhdr_309 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_309_io_clk),
    .io_en(rvclkhdr_309_io_en)
  );
  rvclkhdr rvclkhdr_310 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_310_io_clk),
    .io_en(rvclkhdr_310_io_en)
  );
  rvclkhdr rvclkhdr_311 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_311_io_clk),
    .io_en(rvclkhdr_311_io_en)
  );
  rvclkhdr rvclkhdr_312 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_312_io_clk),
    .io_en(rvclkhdr_312_io_en)
  );
  rvclkhdr rvclkhdr_313 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_313_io_clk),
    .io_en(rvclkhdr_313_io_en)
  );
  rvclkhdr rvclkhdr_314 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_314_io_clk),
    .io_en(rvclkhdr_314_io_en)
  );
  rvclkhdr rvclkhdr_315 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_315_io_clk),
    .io_en(rvclkhdr_315_io_en)
  );
  rvclkhdr rvclkhdr_316 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_316_io_clk),
    .io_en(rvclkhdr_316_io_en)
  );
  rvclkhdr rvclkhdr_317 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_317_io_clk),
    .io_en(rvclkhdr_317_io_en)
  );
  rvclkhdr rvclkhdr_318 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_318_io_clk),
    .io_en(rvclkhdr_318_io_en)
  );
  rvclkhdr rvclkhdr_319 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_319_io_clk),
    .io_en(rvclkhdr_319_io_en)
  );
  rvclkhdr rvclkhdr_320 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_320_io_clk),
    .io_en(rvclkhdr_320_io_en)
  );
  rvclkhdr rvclkhdr_321 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_321_io_clk),
    .io_en(rvclkhdr_321_io_en)
  );
  rvclkhdr rvclkhdr_322 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_322_io_clk),
    .io_en(rvclkhdr_322_io_en)
  );
  rvclkhdr rvclkhdr_323 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_323_io_clk),
    .io_en(rvclkhdr_323_io_en)
  );
  rvclkhdr rvclkhdr_324 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_324_io_clk),
    .io_en(rvclkhdr_324_io_en)
  );
  rvclkhdr rvclkhdr_325 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_325_io_clk),
    .io_en(rvclkhdr_325_io_en)
  );
  rvclkhdr rvclkhdr_326 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_326_io_clk),
    .io_en(rvclkhdr_326_io_en)
  );
  rvclkhdr rvclkhdr_327 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_327_io_clk),
    .io_en(rvclkhdr_327_io_en)
  );
  rvclkhdr rvclkhdr_328 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_328_io_clk),
    .io_en(rvclkhdr_328_io_en)
  );
  rvclkhdr rvclkhdr_329 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_329_io_clk),
    .io_en(rvclkhdr_329_io_en)
  );
  rvclkhdr rvclkhdr_330 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_330_io_clk),
    .io_en(rvclkhdr_330_io_en)
  );
  rvclkhdr rvclkhdr_331 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_331_io_clk),
    .io_en(rvclkhdr_331_io_en)
  );
  rvclkhdr rvclkhdr_332 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_332_io_clk),
    .io_en(rvclkhdr_332_io_en)
  );
  rvclkhdr rvclkhdr_333 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_333_io_clk),
    .io_en(rvclkhdr_333_io_en)
  );
  rvclkhdr rvclkhdr_334 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_334_io_clk),
    .io_en(rvclkhdr_334_io_en)
  );
  rvclkhdr rvclkhdr_335 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_335_io_clk),
    .io_en(rvclkhdr_335_io_en)
  );
  rvclkhdr rvclkhdr_336 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_336_io_clk),
    .io_en(rvclkhdr_336_io_en)
  );
  rvclkhdr rvclkhdr_337 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_337_io_clk),
    .io_en(rvclkhdr_337_io_en)
  );
  rvclkhdr rvclkhdr_338 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_338_io_clk),
    .io_en(rvclkhdr_338_io_en)
  );
  rvclkhdr rvclkhdr_339 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_339_io_clk),
    .io_en(rvclkhdr_339_io_en)
  );
  rvclkhdr rvclkhdr_340 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_340_io_clk),
    .io_en(rvclkhdr_340_io_en)
  );
  rvclkhdr rvclkhdr_341 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_341_io_clk),
    .io_en(rvclkhdr_341_io_en)
  );
  rvclkhdr rvclkhdr_342 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_342_io_clk),
    .io_en(rvclkhdr_342_io_en)
  );
  rvclkhdr rvclkhdr_343 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_343_io_clk),
    .io_en(rvclkhdr_343_io_en)
  );
  rvclkhdr rvclkhdr_344 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_344_io_clk),
    .io_en(rvclkhdr_344_io_en)
  );
  rvclkhdr rvclkhdr_345 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_345_io_clk),
    .io_en(rvclkhdr_345_io_en)
  );
  rvclkhdr rvclkhdr_346 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_346_io_clk),
    .io_en(rvclkhdr_346_io_en)
  );
  rvclkhdr rvclkhdr_347 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_347_io_clk),
    .io_en(rvclkhdr_347_io_en)
  );
  rvclkhdr rvclkhdr_348 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_348_io_clk),
    .io_en(rvclkhdr_348_io_en)
  );
  rvclkhdr rvclkhdr_349 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_349_io_clk),
    .io_en(rvclkhdr_349_io_en)
  );
  rvclkhdr rvclkhdr_350 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_350_io_clk),
    .io_en(rvclkhdr_350_io_en)
  );
  rvclkhdr rvclkhdr_351 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_351_io_clk),
    .io_en(rvclkhdr_351_io_en)
  );
  rvclkhdr rvclkhdr_352 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_352_io_clk),
    .io_en(rvclkhdr_352_io_en)
  );
  rvclkhdr rvclkhdr_353 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_353_io_clk),
    .io_en(rvclkhdr_353_io_en)
  );
  rvclkhdr rvclkhdr_354 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_354_io_clk),
    .io_en(rvclkhdr_354_io_en)
  );
  rvclkhdr rvclkhdr_355 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_355_io_clk),
    .io_en(rvclkhdr_355_io_en)
  );
  rvclkhdr rvclkhdr_356 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_356_io_clk),
    .io_en(rvclkhdr_356_io_en)
  );
  rvclkhdr rvclkhdr_357 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_357_io_clk),
    .io_en(rvclkhdr_357_io_en)
  );
  rvclkhdr rvclkhdr_358 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_358_io_clk),
    .io_en(rvclkhdr_358_io_en)
  );
  rvclkhdr rvclkhdr_359 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_359_io_clk),
    .io_en(rvclkhdr_359_io_en)
  );
  rvclkhdr rvclkhdr_360 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_360_io_clk),
    .io_en(rvclkhdr_360_io_en)
  );
  rvclkhdr rvclkhdr_361 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_361_io_clk),
    .io_en(rvclkhdr_361_io_en)
  );
  rvclkhdr rvclkhdr_362 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_362_io_clk),
    .io_en(rvclkhdr_362_io_en)
  );
  rvclkhdr rvclkhdr_363 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_363_io_clk),
    .io_en(rvclkhdr_363_io_en)
  );
  rvclkhdr rvclkhdr_364 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_364_io_clk),
    .io_en(rvclkhdr_364_io_en)
  );
  rvclkhdr rvclkhdr_365 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_365_io_clk),
    .io_en(rvclkhdr_365_io_en)
  );
  rvclkhdr rvclkhdr_366 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_366_io_clk),
    .io_en(rvclkhdr_366_io_en)
  );
  rvclkhdr rvclkhdr_367 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_367_io_clk),
    .io_en(rvclkhdr_367_io_en)
  );
  rvclkhdr rvclkhdr_368 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_368_io_clk),
    .io_en(rvclkhdr_368_io_en)
  );
  rvclkhdr rvclkhdr_369 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_369_io_clk),
    .io_en(rvclkhdr_369_io_en)
  );
  rvclkhdr rvclkhdr_370 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_370_io_clk),
    .io_en(rvclkhdr_370_io_en)
  );
  rvclkhdr rvclkhdr_371 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_371_io_clk),
    .io_en(rvclkhdr_371_io_en)
  );
  rvclkhdr rvclkhdr_372 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_372_io_clk),
    .io_en(rvclkhdr_372_io_en)
  );
  rvclkhdr rvclkhdr_373 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_373_io_clk),
    .io_en(rvclkhdr_373_io_en)
  );
  rvclkhdr rvclkhdr_374 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_374_io_clk),
    .io_en(rvclkhdr_374_io_en)
  );
  rvclkhdr rvclkhdr_375 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_375_io_clk),
    .io_en(rvclkhdr_375_io_en)
  );
  rvclkhdr rvclkhdr_376 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_376_io_clk),
    .io_en(rvclkhdr_376_io_en)
  );
  rvclkhdr rvclkhdr_377 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_377_io_clk),
    .io_en(rvclkhdr_377_io_en)
  );
  rvclkhdr rvclkhdr_378 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_378_io_clk),
    .io_en(rvclkhdr_378_io_en)
  );
  rvclkhdr rvclkhdr_379 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_379_io_clk),
    .io_en(rvclkhdr_379_io_en)
  );
  rvclkhdr rvclkhdr_380 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_380_io_clk),
    .io_en(rvclkhdr_380_io_en)
  );
  rvclkhdr rvclkhdr_381 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_381_io_clk),
    .io_en(rvclkhdr_381_io_en)
  );
  rvclkhdr rvclkhdr_382 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_382_io_clk),
    .io_en(rvclkhdr_382_io_en)
  );
  rvclkhdr rvclkhdr_383 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_383_io_clk),
    .io_en(rvclkhdr_383_io_en)
  );
  rvclkhdr rvclkhdr_384 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_384_io_clk),
    .io_en(rvclkhdr_384_io_en)
  );
  rvclkhdr rvclkhdr_385 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_385_io_clk),
    .io_en(rvclkhdr_385_io_en)
  );
  rvclkhdr rvclkhdr_386 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_386_io_clk),
    .io_en(rvclkhdr_386_io_en)
  );
  rvclkhdr rvclkhdr_387 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_387_io_clk),
    .io_en(rvclkhdr_387_io_en)
  );
  rvclkhdr rvclkhdr_388 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_388_io_clk),
    .io_en(rvclkhdr_388_io_en)
  );
  rvclkhdr rvclkhdr_389 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_389_io_clk),
    .io_en(rvclkhdr_389_io_en)
  );
  rvclkhdr rvclkhdr_390 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_390_io_clk),
    .io_en(rvclkhdr_390_io_en)
  );
  rvclkhdr rvclkhdr_391 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_391_io_clk),
    .io_en(rvclkhdr_391_io_en)
  );
  rvclkhdr rvclkhdr_392 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_392_io_clk),
    .io_en(rvclkhdr_392_io_en)
  );
  rvclkhdr rvclkhdr_393 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_393_io_clk),
    .io_en(rvclkhdr_393_io_en)
  );
  rvclkhdr rvclkhdr_394 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_394_io_clk),
    .io_en(rvclkhdr_394_io_en)
  );
  rvclkhdr rvclkhdr_395 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_395_io_clk),
    .io_en(rvclkhdr_395_io_en)
  );
  rvclkhdr rvclkhdr_396 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_396_io_clk),
    .io_en(rvclkhdr_396_io_en)
  );
  rvclkhdr rvclkhdr_397 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_397_io_clk),
    .io_en(rvclkhdr_397_io_en)
  );
  rvclkhdr rvclkhdr_398 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_398_io_clk),
    .io_en(rvclkhdr_398_io_en)
  );
  rvclkhdr rvclkhdr_399 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_399_io_clk),
    .io_en(rvclkhdr_399_io_en)
  );
  rvclkhdr rvclkhdr_400 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_400_io_clk),
    .io_en(rvclkhdr_400_io_en)
  );
  rvclkhdr rvclkhdr_401 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_401_io_clk),
    .io_en(rvclkhdr_401_io_en)
  );
  rvclkhdr rvclkhdr_402 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_402_io_clk),
    .io_en(rvclkhdr_402_io_en)
  );
  rvclkhdr rvclkhdr_403 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_403_io_clk),
    .io_en(rvclkhdr_403_io_en)
  );
  rvclkhdr rvclkhdr_404 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_404_io_clk),
    .io_en(rvclkhdr_404_io_en)
  );
  rvclkhdr rvclkhdr_405 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_405_io_clk),
    .io_en(rvclkhdr_405_io_en)
  );
  rvclkhdr rvclkhdr_406 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_406_io_clk),
    .io_en(rvclkhdr_406_io_en)
  );
  rvclkhdr rvclkhdr_407 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_407_io_clk),
    .io_en(rvclkhdr_407_io_en)
  );
  rvclkhdr rvclkhdr_408 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_408_io_clk),
    .io_en(rvclkhdr_408_io_en)
  );
  rvclkhdr rvclkhdr_409 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_409_io_clk),
    .io_en(rvclkhdr_409_io_en)
  );
  rvclkhdr rvclkhdr_410 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_410_io_clk),
    .io_en(rvclkhdr_410_io_en)
  );
  rvclkhdr rvclkhdr_411 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_411_io_clk),
    .io_en(rvclkhdr_411_io_en)
  );
  rvclkhdr rvclkhdr_412 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_412_io_clk),
    .io_en(rvclkhdr_412_io_en)
  );
  rvclkhdr rvclkhdr_413 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_413_io_clk),
    .io_en(rvclkhdr_413_io_en)
  );
  rvclkhdr rvclkhdr_414 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_414_io_clk),
    .io_en(rvclkhdr_414_io_en)
  );
  rvclkhdr rvclkhdr_415 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_415_io_clk),
    .io_en(rvclkhdr_415_io_en)
  );
  rvclkhdr rvclkhdr_416 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_416_io_clk),
    .io_en(rvclkhdr_416_io_en)
  );
  rvclkhdr rvclkhdr_417 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_417_io_clk),
    .io_en(rvclkhdr_417_io_en)
  );
  rvclkhdr rvclkhdr_418 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_418_io_clk),
    .io_en(rvclkhdr_418_io_en)
  );
  rvclkhdr rvclkhdr_419 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_419_io_clk),
    .io_en(rvclkhdr_419_io_en)
  );
  rvclkhdr rvclkhdr_420 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_420_io_clk),
    .io_en(rvclkhdr_420_io_en)
  );
  rvclkhdr rvclkhdr_421 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_421_io_clk),
    .io_en(rvclkhdr_421_io_en)
  );
  rvclkhdr rvclkhdr_422 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_422_io_clk),
    .io_en(rvclkhdr_422_io_en)
  );
  rvclkhdr rvclkhdr_423 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_423_io_clk),
    .io_en(rvclkhdr_423_io_en)
  );
  rvclkhdr rvclkhdr_424 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_424_io_clk),
    .io_en(rvclkhdr_424_io_en)
  );
  rvclkhdr rvclkhdr_425 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_425_io_clk),
    .io_en(rvclkhdr_425_io_en)
  );
  rvclkhdr rvclkhdr_426 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_426_io_clk),
    .io_en(rvclkhdr_426_io_en)
  );
  rvclkhdr rvclkhdr_427 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_427_io_clk),
    .io_en(rvclkhdr_427_io_en)
  );
  rvclkhdr rvclkhdr_428 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_428_io_clk),
    .io_en(rvclkhdr_428_io_en)
  );
  rvclkhdr rvclkhdr_429 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_429_io_clk),
    .io_en(rvclkhdr_429_io_en)
  );
  rvclkhdr rvclkhdr_430 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_430_io_clk),
    .io_en(rvclkhdr_430_io_en)
  );
  rvclkhdr rvclkhdr_431 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_431_io_clk),
    .io_en(rvclkhdr_431_io_en)
  );
  rvclkhdr rvclkhdr_432 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_432_io_clk),
    .io_en(rvclkhdr_432_io_en)
  );
  rvclkhdr rvclkhdr_433 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_433_io_clk),
    .io_en(rvclkhdr_433_io_en)
  );
  rvclkhdr rvclkhdr_434 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_434_io_clk),
    .io_en(rvclkhdr_434_io_en)
  );
  rvclkhdr rvclkhdr_435 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_435_io_clk),
    .io_en(rvclkhdr_435_io_en)
  );
  rvclkhdr rvclkhdr_436 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_436_io_clk),
    .io_en(rvclkhdr_436_io_en)
  );
  rvclkhdr rvclkhdr_437 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_437_io_clk),
    .io_en(rvclkhdr_437_io_en)
  );
  rvclkhdr rvclkhdr_438 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_438_io_clk),
    .io_en(rvclkhdr_438_io_en)
  );
  rvclkhdr rvclkhdr_439 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_439_io_clk),
    .io_en(rvclkhdr_439_io_en)
  );
  rvclkhdr rvclkhdr_440 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_440_io_clk),
    .io_en(rvclkhdr_440_io_en)
  );
  rvclkhdr rvclkhdr_441 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_441_io_clk),
    .io_en(rvclkhdr_441_io_en)
  );
  rvclkhdr rvclkhdr_442 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_442_io_clk),
    .io_en(rvclkhdr_442_io_en)
  );
  rvclkhdr rvclkhdr_443 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_443_io_clk),
    .io_en(rvclkhdr_443_io_en)
  );
  rvclkhdr rvclkhdr_444 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_444_io_clk),
    .io_en(rvclkhdr_444_io_en)
  );
  rvclkhdr rvclkhdr_445 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_445_io_clk),
    .io_en(rvclkhdr_445_io_en)
  );
  rvclkhdr rvclkhdr_446 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_446_io_clk),
    .io_en(rvclkhdr_446_io_en)
  );
  rvclkhdr rvclkhdr_447 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_447_io_clk),
    .io_en(rvclkhdr_447_io_en)
  );
  rvclkhdr rvclkhdr_448 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_448_io_clk),
    .io_en(rvclkhdr_448_io_en)
  );
  rvclkhdr rvclkhdr_449 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_449_io_clk),
    .io_en(rvclkhdr_449_io_en)
  );
  rvclkhdr rvclkhdr_450 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_450_io_clk),
    .io_en(rvclkhdr_450_io_en)
  );
  rvclkhdr rvclkhdr_451 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_451_io_clk),
    .io_en(rvclkhdr_451_io_en)
  );
  rvclkhdr rvclkhdr_452 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_452_io_clk),
    .io_en(rvclkhdr_452_io_en)
  );
  rvclkhdr rvclkhdr_453 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_453_io_clk),
    .io_en(rvclkhdr_453_io_en)
  );
  rvclkhdr rvclkhdr_454 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_454_io_clk),
    .io_en(rvclkhdr_454_io_en)
  );
  rvclkhdr rvclkhdr_455 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_455_io_clk),
    .io_en(rvclkhdr_455_io_en)
  );
  rvclkhdr rvclkhdr_456 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_456_io_clk),
    .io_en(rvclkhdr_456_io_en)
  );
  rvclkhdr rvclkhdr_457 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_457_io_clk),
    .io_en(rvclkhdr_457_io_en)
  );
  rvclkhdr rvclkhdr_458 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_458_io_clk),
    .io_en(rvclkhdr_458_io_en)
  );
  rvclkhdr rvclkhdr_459 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_459_io_clk),
    .io_en(rvclkhdr_459_io_en)
  );
  rvclkhdr rvclkhdr_460 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_460_io_clk),
    .io_en(rvclkhdr_460_io_en)
  );
  rvclkhdr rvclkhdr_461 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_461_io_clk),
    .io_en(rvclkhdr_461_io_en)
  );
  rvclkhdr rvclkhdr_462 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_462_io_clk),
    .io_en(rvclkhdr_462_io_en)
  );
  rvclkhdr rvclkhdr_463 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_463_io_clk),
    .io_en(rvclkhdr_463_io_en)
  );
  rvclkhdr rvclkhdr_464 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_464_io_clk),
    .io_en(rvclkhdr_464_io_en)
  );
  rvclkhdr rvclkhdr_465 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_465_io_clk),
    .io_en(rvclkhdr_465_io_en)
  );
  rvclkhdr rvclkhdr_466 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_466_io_clk),
    .io_en(rvclkhdr_466_io_en)
  );
  rvclkhdr rvclkhdr_467 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_467_io_clk),
    .io_en(rvclkhdr_467_io_en)
  );
  rvclkhdr rvclkhdr_468 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_468_io_clk),
    .io_en(rvclkhdr_468_io_en)
  );
  rvclkhdr rvclkhdr_469 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_469_io_clk),
    .io_en(rvclkhdr_469_io_en)
  );
  rvclkhdr rvclkhdr_470 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_470_io_clk),
    .io_en(rvclkhdr_470_io_en)
  );
  rvclkhdr rvclkhdr_471 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_471_io_clk),
    .io_en(rvclkhdr_471_io_en)
  );
  rvclkhdr rvclkhdr_472 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_472_io_clk),
    .io_en(rvclkhdr_472_io_en)
  );
  rvclkhdr rvclkhdr_473 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_473_io_clk),
    .io_en(rvclkhdr_473_io_en)
  );
  rvclkhdr rvclkhdr_474 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_474_io_clk),
    .io_en(rvclkhdr_474_io_en)
  );
  rvclkhdr rvclkhdr_475 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_475_io_clk),
    .io_en(rvclkhdr_475_io_en)
  );
  rvclkhdr rvclkhdr_476 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_476_io_clk),
    .io_en(rvclkhdr_476_io_en)
  );
  rvclkhdr rvclkhdr_477 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_477_io_clk),
    .io_en(rvclkhdr_477_io_en)
  );
  rvclkhdr rvclkhdr_478 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_478_io_clk),
    .io_en(rvclkhdr_478_io_en)
  );
  rvclkhdr rvclkhdr_479 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_479_io_clk),
    .io_en(rvclkhdr_479_io_en)
  );
  rvclkhdr rvclkhdr_480 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_480_io_clk),
    .io_en(rvclkhdr_480_io_en)
  );
  rvclkhdr rvclkhdr_481 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_481_io_clk),
    .io_en(rvclkhdr_481_io_en)
  );
  rvclkhdr rvclkhdr_482 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_482_io_clk),
    .io_en(rvclkhdr_482_io_en)
  );
  rvclkhdr rvclkhdr_483 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_483_io_clk),
    .io_en(rvclkhdr_483_io_en)
  );
  rvclkhdr rvclkhdr_484 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_484_io_clk),
    .io_en(rvclkhdr_484_io_en)
  );
  rvclkhdr rvclkhdr_485 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_485_io_clk),
    .io_en(rvclkhdr_485_io_en)
  );
  rvclkhdr rvclkhdr_486 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_486_io_clk),
    .io_en(rvclkhdr_486_io_en)
  );
  rvclkhdr rvclkhdr_487 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_487_io_clk),
    .io_en(rvclkhdr_487_io_en)
  );
  rvclkhdr rvclkhdr_488 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_488_io_clk),
    .io_en(rvclkhdr_488_io_en)
  );
  rvclkhdr rvclkhdr_489 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_489_io_clk),
    .io_en(rvclkhdr_489_io_en)
  );
  rvclkhdr rvclkhdr_490 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_490_io_clk),
    .io_en(rvclkhdr_490_io_en)
  );
  rvclkhdr rvclkhdr_491 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_491_io_clk),
    .io_en(rvclkhdr_491_io_en)
  );
  rvclkhdr rvclkhdr_492 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_492_io_clk),
    .io_en(rvclkhdr_492_io_en)
  );
  rvclkhdr rvclkhdr_493 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_493_io_clk),
    .io_en(rvclkhdr_493_io_en)
  );
  rvclkhdr rvclkhdr_494 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_494_io_clk),
    .io_en(rvclkhdr_494_io_en)
  );
  rvclkhdr rvclkhdr_495 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_495_io_clk),
    .io_en(rvclkhdr_495_io_en)
  );
  rvclkhdr rvclkhdr_496 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_496_io_clk),
    .io_en(rvclkhdr_496_io_en)
  );
  rvclkhdr rvclkhdr_497 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_497_io_clk),
    .io_en(rvclkhdr_497_io_en)
  );
  rvclkhdr rvclkhdr_498 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_498_io_clk),
    .io_en(rvclkhdr_498_io_en)
  );
  rvclkhdr rvclkhdr_499 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_499_io_clk),
    .io_en(rvclkhdr_499_io_en)
  );
  rvclkhdr rvclkhdr_500 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_500_io_clk),
    .io_en(rvclkhdr_500_io_en)
  );
  rvclkhdr rvclkhdr_501 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_501_io_clk),
    .io_en(rvclkhdr_501_io_en)
  );
  rvclkhdr rvclkhdr_502 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_502_io_clk),
    .io_en(rvclkhdr_502_io_en)
  );
  rvclkhdr rvclkhdr_503 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_503_io_clk),
    .io_en(rvclkhdr_503_io_en)
  );
  rvclkhdr rvclkhdr_504 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_504_io_clk),
    .io_en(rvclkhdr_504_io_en)
  );
  rvclkhdr rvclkhdr_505 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_505_io_clk),
    .io_en(rvclkhdr_505_io_en)
  );
  rvclkhdr rvclkhdr_506 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_506_io_clk),
    .io_en(rvclkhdr_506_io_en)
  );
  rvclkhdr rvclkhdr_507 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_507_io_clk),
    .io_en(rvclkhdr_507_io_en)
  );
  rvclkhdr rvclkhdr_508 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_508_io_clk),
    .io_en(rvclkhdr_508_io_en)
  );
  rvclkhdr rvclkhdr_509 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_509_io_clk),
    .io_en(rvclkhdr_509_io_en)
  );
  rvclkhdr rvclkhdr_510 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_510_io_clk),
    .io_en(rvclkhdr_510_io_en)
  );
  rvclkhdr rvclkhdr_511 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_511_io_clk),
    .io_en(rvclkhdr_511_io_en)
  );
  rvclkhdr rvclkhdr_512 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_512_io_clk),
    .io_en(rvclkhdr_512_io_en)
  );
  rvclkhdr rvclkhdr_513 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_513_io_clk),
    .io_en(rvclkhdr_513_io_en)
  );
  rvclkhdr rvclkhdr_514 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_514_io_clk),
    .io_en(rvclkhdr_514_io_en)
  );
  rvclkhdr rvclkhdr_515 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_515_io_clk),
    .io_en(rvclkhdr_515_io_en)
  );
  rvclkhdr rvclkhdr_516 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_516_io_clk),
    .io_en(rvclkhdr_516_io_en)
  );
  rvclkhdr rvclkhdr_517 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_517_io_clk),
    .io_en(rvclkhdr_517_io_en)
  );
  rvclkhdr rvclkhdr_518 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_518_io_clk),
    .io_en(rvclkhdr_518_io_en)
  );
  rvclkhdr rvclkhdr_519 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_519_io_clk),
    .io_en(rvclkhdr_519_io_en)
  );
  rvclkhdr rvclkhdr_520 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_520_io_clk),
    .io_en(rvclkhdr_520_io_en)
  );
  rvclkhdr rvclkhdr_521 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_521_io_clk),
    .io_en(rvclkhdr_521_io_en)
  );
  rvclkhdr rvclkhdr_522 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_522_io_clk),
    .io_en(rvclkhdr_522_io_en)
  );
  rvclkhdr rvclkhdr_523 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_523_io_clk),
    .io_en(rvclkhdr_523_io_en)
  );
  rvclkhdr rvclkhdr_524 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_524_io_clk),
    .io_en(rvclkhdr_524_io_en)
  );
  rvclkhdr rvclkhdr_525 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_525_io_clk),
    .io_en(rvclkhdr_525_io_en)
  );
  rvclkhdr rvclkhdr_526 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_526_io_clk),
    .io_en(rvclkhdr_526_io_en)
  );
  rvclkhdr rvclkhdr_527 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_527_io_clk),
    .io_en(rvclkhdr_527_io_en)
  );
  rvclkhdr rvclkhdr_528 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_528_io_clk),
    .io_en(rvclkhdr_528_io_en)
  );
  rvclkhdr rvclkhdr_529 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_529_io_clk),
    .io_en(rvclkhdr_529_io_en)
  );
  rvclkhdr rvclkhdr_530 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_530_io_clk),
    .io_en(rvclkhdr_530_io_en)
  );
  rvclkhdr rvclkhdr_531 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_531_io_clk),
    .io_en(rvclkhdr_531_io_en)
  );
  rvclkhdr rvclkhdr_532 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_532_io_clk),
    .io_en(rvclkhdr_532_io_en)
  );
  rvclkhdr rvclkhdr_533 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_533_io_clk),
    .io_en(rvclkhdr_533_io_en)
  );
  rvclkhdr rvclkhdr_534 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_534_io_clk),
    .io_en(rvclkhdr_534_io_en)
  );
  rvclkhdr rvclkhdr_535 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_535_io_clk),
    .io_en(rvclkhdr_535_io_en)
  );
  rvclkhdr rvclkhdr_536 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_536_io_clk),
    .io_en(rvclkhdr_536_io_en)
  );
  rvclkhdr rvclkhdr_537 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_537_io_clk),
    .io_en(rvclkhdr_537_io_en)
  );
  rvclkhdr rvclkhdr_538 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_538_io_clk),
    .io_en(rvclkhdr_538_io_en)
  );
  rvclkhdr rvclkhdr_539 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_539_io_clk),
    .io_en(rvclkhdr_539_io_en)
  );
  rvclkhdr rvclkhdr_540 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_540_io_clk),
    .io_en(rvclkhdr_540_io_en)
  );
  rvclkhdr rvclkhdr_541 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_541_io_clk),
    .io_en(rvclkhdr_541_io_en)
  );
  rvclkhdr rvclkhdr_542 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_542_io_clk),
    .io_en(rvclkhdr_542_io_en)
  );
  rvclkhdr rvclkhdr_543 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_543_io_clk),
    .io_en(rvclkhdr_543_io_en)
  );
  rvclkhdr rvclkhdr_544 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_544_io_clk),
    .io_en(rvclkhdr_544_io_en)
  );
  rvclkhdr rvclkhdr_545 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_545_io_clk),
    .io_en(rvclkhdr_545_io_en)
  );
  rvclkhdr rvclkhdr_546 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_546_io_clk),
    .io_en(rvclkhdr_546_io_en)
  );
  rvclkhdr rvclkhdr_547 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_547_io_clk),
    .io_en(rvclkhdr_547_io_en)
  );
  rvclkhdr rvclkhdr_548 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_548_io_clk),
    .io_en(rvclkhdr_548_io_en)
  );
  rvclkhdr rvclkhdr_549 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_549_io_clk),
    .io_en(rvclkhdr_549_io_en)
  );
  rvclkhdr rvclkhdr_550 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_550_io_clk),
    .io_en(rvclkhdr_550_io_en)
  );
  rvclkhdr rvclkhdr_551 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_551_io_clk),
    .io_en(rvclkhdr_551_io_en)
  );
  rvclkhdr rvclkhdr_552 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_552_io_clk),
    .io_en(rvclkhdr_552_io_en)
  );
  assign io_ifu_bp_hit_taken_f = _T_257 & _T_258; // @[ifu_bp_ctl.scala 277:25]
  assign io_ifu_bp_btb_target_f = _T_469 | _T_479; // @[ifu_bp_ctl.scala 374:26]
  assign io_ifu_bp_inst_mask_f = _T_294 | _T_295; // @[ifu_bp_ctl.scala 302:25]
  assign io_ifu_bp_fghr_f = fghr; // @[ifu_bp_ctl.scala 345:20]
  assign io_ifu_bp_way_f = tag_match_vway1_expanded_f | _T_169; // @[ifu_bp_ctl.scala 254:19]
  assign io_ifu_bp_ret_f = {_T_314,_T_320}; // @[ifu_bp_ctl.scala 351:19]
  assign io_ifu_bp_hist1_f = bht_force_taken_f | _T_299; // @[ifu_bp_ctl.scala 346:21]
  assign io_ifu_bp_hist0_f = {bht_vbank1_rd_data_f[0],bht_vbank0_rd_data_f[0]}; // @[ifu_bp_ctl.scala 347:21]
  assign io_ifu_bp_pc4_f = {_T_305,_T_308}; // @[ifu_bp_ctl.scala 348:19]
  assign io_ifu_bp_valid_f = bht_valid_f & _T_379; // @[ifu_bp_ctl.scala 350:21]
  assign io_ifu_bp_poffset_f = btb_sel_data_f[15:4]; // @[ifu_bp_ctl.scala 362:23]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_io_en = io_ifc_fetch_req_f | exu_mp_valid; // @[lib.scala 412:17]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_1_io_en = ~rs_hold; // @[lib.scala 412:17]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_2_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_3_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_4_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_5_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_6_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_7_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_8_io_en = _T_520 & io_ifu_bp_hit_taken_f; // @[lib.scala 412:17]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_9_io_en = _T_642 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_10_io_en = _T_646 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_11_io_en = _T_650 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_12_io_en = _T_654 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_13_io_en = _T_658 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_14_io_en = _T_662 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_15_io_en = _T_666 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_16_io_en = _T_670 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_17_io_en = _T_674 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_18_io_en = _T_678 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_19_io_en = _T_682 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_20_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_20_io_en = _T_686 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_21_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_21_io_en = _T_690 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_22_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_22_io_en = _T_694 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_23_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_23_io_en = _T_698 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_24_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_24_io_en = _T_702 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_25_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_25_io_en = _T_706 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_26_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_26_io_en = _T_710 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_27_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_27_io_en = _T_714 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_28_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_28_io_en = _T_718 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_29_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_29_io_en = _T_722 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_30_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_30_io_en = _T_726 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_31_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_31_io_en = _T_730 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_32_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_32_io_en = _T_734 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_33_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_33_io_en = _T_738 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_34_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_34_io_en = _T_742 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_35_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_35_io_en = _T_746 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_36_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_36_io_en = _T_750 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_37_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_37_io_en = _T_754 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_38_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_38_io_en = _T_758 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_39_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_39_io_en = _T_762 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_40_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_40_io_en = _T_766 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_41_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_41_io_en = _T_770 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_42_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_42_io_en = _T_774 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_43_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_43_io_en = _T_778 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_44_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_44_io_en = _T_782 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_45_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_45_io_en = _T_786 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_46_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_46_io_en = _T_790 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_47_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_47_io_en = _T_794 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_48_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_48_io_en = _T_798 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_49_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_49_io_en = _T_802 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_50_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_50_io_en = _T_806 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_51_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_51_io_en = _T_810 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_52_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_52_io_en = _T_814 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_53_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_53_io_en = _T_818 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_54_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_54_io_en = _T_822 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_55_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_55_io_en = _T_826 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_56_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_56_io_en = _T_830 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_57_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_57_io_en = _T_834 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_58_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_58_io_en = _T_838 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_59_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_59_io_en = _T_842 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_60_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_60_io_en = _T_846 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_61_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_61_io_en = _T_850 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_62_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_62_io_en = _T_854 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_63_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_63_io_en = _T_858 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_64_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_64_io_en = _T_862 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_65_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_65_io_en = _T_866 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_66_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_66_io_en = _T_870 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_67_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_67_io_en = _T_874 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_68_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_68_io_en = _T_878 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_69_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_69_io_en = _T_882 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_70_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_70_io_en = _T_886 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_71_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_71_io_en = _T_890 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_72_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_72_io_en = _T_894 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_73_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_73_io_en = _T_898 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_74_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_74_io_en = _T_902 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_75_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_75_io_en = _T_906 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_76_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_76_io_en = _T_910 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_77_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_77_io_en = _T_914 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_78_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_78_io_en = _T_918 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_79_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_79_io_en = _T_922 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_80_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_80_io_en = _T_926 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_81_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_81_io_en = _T_930 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_82_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_82_io_en = _T_934 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_83_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_83_io_en = _T_938 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_84_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_84_io_en = _T_942 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_85_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_85_io_en = _T_946 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_86_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_86_io_en = _T_950 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_87_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_87_io_en = _T_954 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_88_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_88_io_en = _T_958 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_89_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_89_io_en = _T_962 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_90_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_90_io_en = _T_966 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_91_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_91_io_en = _T_970 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_92_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_92_io_en = _T_974 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_93_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_93_io_en = _T_978 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_94_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_94_io_en = _T_982 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_95_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_95_io_en = _T_986 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_96_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_96_io_en = _T_990 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_97_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_97_io_en = _T_994 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_98_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_98_io_en = _T_998 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_99_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_99_io_en = _T_1002 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_100_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_100_io_en = _T_1006 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_101_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_101_io_en = _T_1010 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_102_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_102_io_en = _T_1014 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_103_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_103_io_en = _T_1018 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_104_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_104_io_en = _T_1022 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_105_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_105_io_en = _T_1026 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_106_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_106_io_en = _T_1030 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_107_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_107_io_en = _T_1034 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_108_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_108_io_en = _T_1038 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_109_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_109_io_en = _T_1042 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_110_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_110_io_en = _T_1046 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_111_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_111_io_en = _T_1050 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_112_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_112_io_en = _T_1054 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_113_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_113_io_en = _T_1058 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_114_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_114_io_en = _T_1062 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_115_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_115_io_en = _T_1066 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_116_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_116_io_en = _T_1070 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_117_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_117_io_en = _T_1074 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_118_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_118_io_en = _T_1078 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_119_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_119_io_en = _T_1082 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_120_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_120_io_en = _T_1086 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_121_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_121_io_en = _T_1090 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_122_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_122_io_en = _T_1094 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_123_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_123_io_en = _T_1098 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_124_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_124_io_en = _T_1102 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_125_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_125_io_en = _T_1106 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_126_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_126_io_en = _T_1110 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_127_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_127_io_en = _T_1114 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_128_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_128_io_en = _T_1118 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_129_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_129_io_en = _T_1122 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_130_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_130_io_en = _T_1126 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_131_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_131_io_en = _T_1130 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_132_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_132_io_en = _T_1134 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_133_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_133_io_en = _T_1138 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_134_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_134_io_en = _T_1142 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_135_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_135_io_en = _T_1146 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_136_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_136_io_en = _T_1150 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_137_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_137_io_en = _T_1154 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_138_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_138_io_en = _T_1158 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_139_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_139_io_en = _T_1162 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_140_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_140_io_en = _T_1166 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_141_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_141_io_en = _T_1170 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_142_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_142_io_en = _T_1174 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_143_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_143_io_en = _T_1178 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_144_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_144_io_en = _T_1182 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_145_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_145_io_en = _T_1186 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_146_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_146_io_en = _T_1190 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_147_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_147_io_en = _T_1194 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_148_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_148_io_en = _T_1198 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_149_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_149_io_en = _T_1202 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_150_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_150_io_en = _T_1206 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_151_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_151_io_en = _T_1210 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_152_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_152_io_en = _T_1214 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_153_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_153_io_en = _T_1218 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_154_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_154_io_en = _T_1222 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_155_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_155_io_en = _T_1226 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_156_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_156_io_en = _T_1230 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_157_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_157_io_en = _T_1234 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_158_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_158_io_en = _T_1238 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_159_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_159_io_en = _T_1242 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_160_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_160_io_en = _T_1246 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_161_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_161_io_en = _T_1250 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_162_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_162_io_en = _T_1254 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_163_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_163_io_en = _T_1258 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_164_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_164_io_en = _T_1262 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_165_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_165_io_en = _T_1266 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_166_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_166_io_en = _T_1270 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_167_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_167_io_en = _T_1274 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_168_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_168_io_en = _T_1278 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_169_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_169_io_en = _T_1282 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_170_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_170_io_en = _T_1286 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_171_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_171_io_en = _T_1290 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_172_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_172_io_en = _T_1294 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_173_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_173_io_en = _T_1298 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_174_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_174_io_en = _T_1302 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_175_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_175_io_en = _T_1306 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_176_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_176_io_en = _T_1310 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_177_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_177_io_en = _T_1314 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_178_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_178_io_en = _T_1318 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_179_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_179_io_en = _T_1322 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_180_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_180_io_en = _T_1326 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_181_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_181_io_en = _T_1330 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_182_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_182_io_en = _T_1334 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_183_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_183_io_en = _T_1338 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_184_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_184_io_en = _T_1342 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_185_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_185_io_en = _T_1346 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_186_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_186_io_en = _T_1350 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_187_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_187_io_en = _T_1354 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_188_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_188_io_en = _T_1358 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_189_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_189_io_en = _T_1362 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_190_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_190_io_en = _T_1366 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_191_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_191_io_en = _T_1370 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_192_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_192_io_en = _T_1374 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_193_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_193_io_en = _T_1378 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_194_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_194_io_en = _T_1382 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_195_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_195_io_en = _T_1386 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_196_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_196_io_en = _T_1390 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_197_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_197_io_en = _T_1394 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_198_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_198_io_en = _T_1398 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_199_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_199_io_en = _T_1402 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_200_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_200_io_en = _T_1406 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_201_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_201_io_en = _T_1410 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_202_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_202_io_en = _T_1414 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_203_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_203_io_en = _T_1418 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_204_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_204_io_en = _T_1422 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_205_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_205_io_en = _T_1426 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_206_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_206_io_en = _T_1430 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_207_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_207_io_en = _T_1434 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_208_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_208_io_en = _T_1438 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_209_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_209_io_en = _T_1442 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_210_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_210_io_en = _T_1446 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_211_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_211_io_en = _T_1450 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_212_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_212_io_en = _T_1454 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_213_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_213_io_en = _T_1458 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_214_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_214_io_en = _T_1462 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_215_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_215_io_en = _T_1466 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_216_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_216_io_en = _T_1470 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_217_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_217_io_en = _T_1474 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_218_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_218_io_en = _T_1478 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_219_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_219_io_en = _T_1482 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_220_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_220_io_en = _T_1486 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_221_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_221_io_en = _T_1490 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_222_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_222_io_en = _T_1494 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_223_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_223_io_en = _T_1498 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_224_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_224_io_en = _T_1502 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_225_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_225_io_en = _T_1506 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_226_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_226_io_en = _T_1510 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_227_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_227_io_en = _T_1514 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_228_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_228_io_en = _T_1518 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_229_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_229_io_en = _T_1522 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_230_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_230_io_en = _T_1526 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_231_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_231_io_en = _T_1530 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_232_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_232_io_en = _T_1534 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_233_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_233_io_en = _T_1538 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_234_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_234_io_en = _T_1542 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_235_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_235_io_en = _T_1546 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_236_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_236_io_en = _T_1550 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_237_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_237_io_en = _T_1554 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_238_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_238_io_en = _T_1558 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_239_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_239_io_en = _T_1562 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_240_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_240_io_en = _T_1566 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_241_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_241_io_en = _T_1570 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_242_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_242_io_en = _T_1574 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_243_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_243_io_en = _T_1578 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_244_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_244_io_en = _T_1582 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_245_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_245_io_en = _T_1586 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_246_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_246_io_en = _T_1590 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_247_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_247_io_en = _T_1594 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_248_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_248_io_en = _T_1598 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_249_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_249_io_en = _T_1602 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_250_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_250_io_en = _T_1606 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_251_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_251_io_en = _T_1610 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_252_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_252_io_en = _T_1614 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_253_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_253_io_en = _T_1618 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_254_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_254_io_en = _T_1622 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_255_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_255_io_en = _T_1626 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_256_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_256_io_en = _T_1630 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_257_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_257_io_en = _T_1634 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_258_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_258_io_en = _T_1638 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_259_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_259_io_en = _T_1642 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_260_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_260_io_en = _T_1646 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_261_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_261_io_en = _T_1650 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_262_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_262_io_en = _T_1654 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_263_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_263_io_en = _T_1658 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_264_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_264_io_en = _T_1662 & _T_620; // @[lib.scala 412:17]
  assign rvclkhdr_265_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_265_io_en = _T_642 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_266_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_266_io_en = _T_646 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_267_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_267_io_en = _T_650 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_268_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_268_io_en = _T_654 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_269_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_269_io_en = _T_658 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_270_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_270_io_en = _T_662 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_271_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_271_io_en = _T_666 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_272_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_272_io_en = _T_670 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_273_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_273_io_en = _T_674 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_274_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_274_io_en = _T_678 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_275_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_275_io_en = _T_682 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_276_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_276_io_en = _T_686 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_277_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_277_io_en = _T_690 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_278_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_278_io_en = _T_694 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_279_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_279_io_en = _T_698 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_280_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_280_io_en = _T_702 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_281_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_281_io_en = _T_706 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_282_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_282_io_en = _T_710 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_283_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_283_io_en = _T_714 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_284_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_284_io_en = _T_718 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_285_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_285_io_en = _T_722 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_286_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_286_io_en = _T_726 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_287_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_287_io_en = _T_730 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_288_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_288_io_en = _T_734 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_289_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_289_io_en = _T_738 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_290_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_290_io_en = _T_742 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_291_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_291_io_en = _T_746 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_292_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_292_io_en = _T_750 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_293_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_293_io_en = _T_754 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_294_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_294_io_en = _T_758 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_295_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_295_io_en = _T_762 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_296_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_296_io_en = _T_766 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_297_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_297_io_en = _T_770 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_298_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_298_io_en = _T_774 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_299_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_299_io_en = _T_778 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_300_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_300_io_en = _T_782 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_301_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_301_io_en = _T_786 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_302_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_302_io_en = _T_790 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_303_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_303_io_en = _T_794 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_304_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_304_io_en = _T_798 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_305_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_305_io_en = _T_802 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_306_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_306_io_en = _T_806 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_307_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_307_io_en = _T_810 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_308_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_308_io_en = _T_814 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_309_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_309_io_en = _T_818 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_310_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_310_io_en = _T_822 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_311_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_311_io_en = _T_826 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_312_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_312_io_en = _T_830 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_313_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_313_io_en = _T_834 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_314_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_314_io_en = _T_838 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_315_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_315_io_en = _T_842 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_316_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_316_io_en = _T_846 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_317_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_317_io_en = _T_850 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_318_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_318_io_en = _T_854 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_319_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_319_io_en = _T_858 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_320_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_320_io_en = _T_862 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_321_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_321_io_en = _T_866 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_322_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_322_io_en = _T_870 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_323_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_323_io_en = _T_874 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_324_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_324_io_en = _T_878 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_325_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_325_io_en = _T_882 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_326_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_326_io_en = _T_886 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_327_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_327_io_en = _T_890 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_328_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_328_io_en = _T_894 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_329_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_329_io_en = _T_898 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_330_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_330_io_en = _T_902 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_331_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_331_io_en = _T_906 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_332_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_332_io_en = _T_910 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_333_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_333_io_en = _T_914 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_334_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_334_io_en = _T_918 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_335_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_335_io_en = _T_922 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_336_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_336_io_en = _T_926 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_337_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_337_io_en = _T_930 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_338_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_338_io_en = _T_934 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_339_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_339_io_en = _T_938 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_340_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_340_io_en = _T_942 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_341_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_341_io_en = _T_946 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_342_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_342_io_en = _T_950 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_343_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_343_io_en = _T_954 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_344_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_344_io_en = _T_958 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_345_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_345_io_en = _T_962 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_346_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_346_io_en = _T_966 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_347_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_347_io_en = _T_970 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_348_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_348_io_en = _T_974 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_349_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_349_io_en = _T_978 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_350_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_350_io_en = _T_982 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_351_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_351_io_en = _T_986 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_352_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_352_io_en = _T_990 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_353_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_353_io_en = _T_994 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_354_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_354_io_en = _T_998 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_355_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_355_io_en = _T_1002 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_356_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_356_io_en = _T_1006 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_357_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_357_io_en = _T_1010 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_358_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_358_io_en = _T_1014 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_359_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_359_io_en = _T_1018 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_360_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_360_io_en = _T_1022 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_361_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_361_io_en = _T_1026 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_362_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_362_io_en = _T_1030 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_363_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_363_io_en = _T_1034 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_364_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_364_io_en = _T_1038 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_365_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_365_io_en = _T_1042 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_366_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_366_io_en = _T_1046 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_367_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_367_io_en = _T_1050 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_368_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_368_io_en = _T_1054 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_369_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_369_io_en = _T_1058 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_370_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_370_io_en = _T_1062 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_371_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_371_io_en = _T_1066 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_372_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_372_io_en = _T_1070 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_373_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_373_io_en = _T_1074 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_374_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_374_io_en = _T_1078 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_375_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_375_io_en = _T_1082 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_376_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_376_io_en = _T_1086 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_377_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_377_io_en = _T_1090 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_378_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_378_io_en = _T_1094 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_379_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_379_io_en = _T_1098 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_380_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_380_io_en = _T_1102 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_381_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_381_io_en = _T_1106 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_382_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_382_io_en = _T_1110 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_383_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_383_io_en = _T_1114 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_384_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_384_io_en = _T_1118 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_385_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_385_io_en = _T_1122 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_386_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_386_io_en = _T_1126 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_387_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_387_io_en = _T_1130 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_388_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_388_io_en = _T_1134 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_389_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_389_io_en = _T_1138 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_390_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_390_io_en = _T_1142 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_391_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_391_io_en = _T_1146 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_392_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_392_io_en = _T_1150 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_393_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_393_io_en = _T_1154 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_394_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_394_io_en = _T_1158 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_395_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_395_io_en = _T_1162 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_396_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_396_io_en = _T_1166 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_397_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_397_io_en = _T_1170 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_398_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_398_io_en = _T_1174 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_399_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_399_io_en = _T_1178 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_400_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_400_io_en = _T_1182 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_401_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_401_io_en = _T_1186 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_402_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_402_io_en = _T_1190 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_403_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_403_io_en = _T_1194 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_404_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_404_io_en = _T_1198 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_405_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_405_io_en = _T_1202 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_406_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_406_io_en = _T_1206 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_407_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_407_io_en = _T_1210 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_408_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_408_io_en = _T_1214 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_409_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_409_io_en = _T_1218 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_410_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_410_io_en = _T_1222 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_411_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_411_io_en = _T_1226 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_412_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_412_io_en = _T_1230 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_413_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_413_io_en = _T_1234 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_414_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_414_io_en = _T_1238 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_415_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_415_io_en = _T_1242 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_416_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_416_io_en = _T_1246 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_417_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_417_io_en = _T_1250 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_418_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_418_io_en = _T_1254 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_419_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_419_io_en = _T_1258 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_420_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_420_io_en = _T_1262 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_421_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_421_io_en = _T_1266 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_422_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_422_io_en = _T_1270 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_423_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_423_io_en = _T_1274 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_424_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_424_io_en = _T_1278 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_425_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_425_io_en = _T_1282 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_426_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_426_io_en = _T_1286 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_427_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_427_io_en = _T_1290 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_428_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_428_io_en = _T_1294 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_429_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_429_io_en = _T_1298 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_430_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_430_io_en = _T_1302 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_431_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_431_io_en = _T_1306 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_432_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_432_io_en = _T_1310 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_433_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_433_io_en = _T_1314 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_434_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_434_io_en = _T_1318 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_435_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_435_io_en = _T_1322 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_436_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_436_io_en = _T_1326 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_437_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_437_io_en = _T_1330 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_438_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_438_io_en = _T_1334 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_439_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_439_io_en = _T_1338 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_440_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_440_io_en = _T_1342 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_441_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_441_io_en = _T_1346 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_442_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_442_io_en = _T_1350 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_443_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_443_io_en = _T_1354 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_444_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_444_io_en = _T_1358 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_445_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_445_io_en = _T_1362 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_446_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_446_io_en = _T_1366 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_447_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_447_io_en = _T_1370 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_448_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_448_io_en = _T_1374 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_449_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_449_io_en = _T_1378 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_450_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_450_io_en = _T_1382 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_451_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_451_io_en = _T_1386 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_452_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_452_io_en = _T_1390 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_453_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_453_io_en = _T_1394 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_454_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_454_io_en = _T_1398 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_455_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_455_io_en = _T_1402 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_456_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_456_io_en = _T_1406 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_457_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_457_io_en = _T_1410 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_458_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_458_io_en = _T_1414 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_459_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_459_io_en = _T_1418 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_460_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_460_io_en = _T_1422 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_461_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_461_io_en = _T_1426 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_462_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_462_io_en = _T_1430 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_463_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_463_io_en = _T_1434 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_464_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_464_io_en = _T_1438 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_465_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_465_io_en = _T_1442 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_466_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_466_io_en = _T_1446 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_467_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_467_io_en = _T_1450 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_468_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_468_io_en = _T_1454 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_469_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_469_io_en = _T_1458 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_470_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_470_io_en = _T_1462 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_471_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_471_io_en = _T_1466 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_472_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_472_io_en = _T_1470 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_473_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_473_io_en = _T_1474 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_474_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_474_io_en = _T_1478 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_475_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_475_io_en = _T_1482 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_476_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_476_io_en = _T_1486 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_477_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_477_io_en = _T_1490 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_478_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_478_io_en = _T_1494 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_479_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_479_io_en = _T_1498 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_480_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_480_io_en = _T_1502 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_481_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_481_io_en = _T_1506 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_482_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_482_io_en = _T_1510 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_483_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_483_io_en = _T_1514 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_484_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_484_io_en = _T_1518 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_485_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_485_io_en = _T_1522 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_486_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_486_io_en = _T_1526 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_487_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_487_io_en = _T_1530 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_488_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_488_io_en = _T_1534 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_489_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_489_io_en = _T_1538 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_490_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_490_io_en = _T_1542 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_491_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_491_io_en = _T_1546 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_492_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_492_io_en = _T_1550 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_493_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_493_io_en = _T_1554 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_494_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_494_io_en = _T_1558 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_495_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_495_io_en = _T_1562 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_496_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_496_io_en = _T_1566 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_497_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_497_io_en = _T_1570 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_498_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_498_io_en = _T_1574 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_499_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_499_io_en = _T_1578 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_500_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_500_io_en = _T_1582 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_501_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_501_io_en = _T_1586 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_502_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_502_io_en = _T_1590 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_503_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_503_io_en = _T_1594 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_504_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_504_io_en = _T_1598 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_505_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_505_io_en = _T_1602 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_506_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_506_io_en = _T_1606 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_507_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_507_io_en = _T_1610 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_508_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_508_io_en = _T_1614 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_509_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_509_io_en = _T_1618 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_510_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_510_io_en = _T_1622 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_511_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_511_io_en = _T_1626 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_512_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_512_io_en = _T_1630 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_513_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_513_io_en = _T_1634 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_514_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_514_io_en = _T_1638 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_515_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_515_io_en = _T_1642 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_516_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_516_io_en = _T_1646 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_517_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_517_io_en = _T_1650 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_518_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_518_io_en = _T_1654 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_519_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_519_io_en = _T_1658 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_520_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_520_io_en = _T_1662 & _T_625; // @[lib.scala 412:17]
  assign rvclkhdr_521_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_521_io_en = _T_6790 | _T_6795; // @[lib.scala 345:16]
  assign rvclkhdr_522_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_522_io_en = _T_6801 | _T_6806; // @[lib.scala 345:16]
  assign rvclkhdr_523_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_523_io_en = _T_6812 | _T_6817; // @[lib.scala 345:16]
  assign rvclkhdr_524_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_524_io_en = _T_6823 | _T_6828; // @[lib.scala 345:16]
  assign rvclkhdr_525_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_525_io_en = _T_6834 | _T_6839; // @[lib.scala 345:16]
  assign rvclkhdr_526_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_526_io_en = _T_6845 | _T_6850; // @[lib.scala 345:16]
  assign rvclkhdr_527_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_527_io_en = _T_6856 | _T_6861; // @[lib.scala 345:16]
  assign rvclkhdr_528_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_528_io_en = _T_6867 | _T_6872; // @[lib.scala 345:16]
  assign rvclkhdr_529_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_529_io_en = _T_6878 | _T_6883; // @[lib.scala 345:16]
  assign rvclkhdr_530_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_530_io_en = _T_6889 | _T_6894; // @[lib.scala 345:16]
  assign rvclkhdr_531_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_531_io_en = _T_6900 | _T_6905; // @[lib.scala 345:16]
  assign rvclkhdr_532_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_532_io_en = _T_6911 | _T_6916; // @[lib.scala 345:16]
  assign rvclkhdr_533_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_533_io_en = _T_6922 | _T_6927; // @[lib.scala 345:16]
  assign rvclkhdr_534_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_534_io_en = _T_6933 | _T_6938; // @[lib.scala 345:16]
  assign rvclkhdr_535_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_535_io_en = _T_6944 | _T_6949; // @[lib.scala 345:16]
  assign rvclkhdr_536_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_536_io_en = _T_6955 | _T_6960; // @[lib.scala 345:16]
  assign rvclkhdr_537_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_537_io_en = _T_6966 | _T_6971; // @[lib.scala 345:16]
  assign rvclkhdr_538_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_538_io_en = _T_6977 | _T_6982; // @[lib.scala 345:16]
  assign rvclkhdr_539_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_539_io_en = _T_6988 | _T_6993; // @[lib.scala 345:16]
  assign rvclkhdr_540_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_540_io_en = _T_6999 | _T_7004; // @[lib.scala 345:16]
  assign rvclkhdr_541_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_541_io_en = _T_7010 | _T_7015; // @[lib.scala 345:16]
  assign rvclkhdr_542_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_542_io_en = _T_7021 | _T_7026; // @[lib.scala 345:16]
  assign rvclkhdr_543_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_543_io_en = _T_7032 | _T_7037; // @[lib.scala 345:16]
  assign rvclkhdr_544_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_544_io_en = _T_7043 | _T_7048; // @[lib.scala 345:16]
  assign rvclkhdr_545_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_545_io_en = _T_7054 | _T_7059; // @[lib.scala 345:16]
  assign rvclkhdr_546_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_546_io_en = _T_7065 | _T_7070; // @[lib.scala 345:16]
  assign rvclkhdr_547_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_547_io_en = _T_7076 | _T_7081; // @[lib.scala 345:16]
  assign rvclkhdr_548_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_548_io_en = _T_7087 | _T_7092; // @[lib.scala 345:16]
  assign rvclkhdr_549_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_549_io_en = _T_7098 | _T_7103; // @[lib.scala 345:16]
  assign rvclkhdr_550_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_550_io_en = _T_7109 | _T_7114; // @[lib.scala 345:16]
  assign rvclkhdr_551_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_551_io_en = _T_7120 | _T_7125; // @[lib.scala 345:16]
  assign rvclkhdr_552_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_552_io_en = _T_7131 | _T_7136; // @[lib.scala 345:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  leak_one_f_d1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_645 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  _T_649 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  _T_653 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  _T_657 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  _T_661 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  _T_665 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  _T_669 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  _T_673 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  _T_677 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  _T_681 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  _T_685 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  _T_689 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  _T_693 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  _T_697 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  _T_701 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  _T_705 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  _T_709 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  _T_713 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  _T_717 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  _T_721 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  _T_725 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  _T_729 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  _T_733 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  _T_737 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  _T_741 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  _T_745 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  _T_749 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  _T_753 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  _T_757 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  _T_761 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  _T_765 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  _T_769 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  _T_773 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  _T_777 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  _T_781 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  _T_785 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  _T_789 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  _T_793 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  _T_797 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  _T_801 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  _T_805 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  _T_809 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  _T_813 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  _T_817 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  _T_821 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  _T_825 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  _T_829 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  _T_833 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  _T_837 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  _T_841 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  _T_845 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  _T_849 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  _T_853 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  _T_857 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  _T_861 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  _T_865 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  _T_869 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  _T_873 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  _T_877 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  _T_881 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  _T_885 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  _T_889 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  _T_893 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  _T_897 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  _T_901 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  _T_905 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  _T_909 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  _T_913 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  _T_917 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  _T_921 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  _T_925 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  _T_929 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  _T_933 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  _T_937 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  _T_941 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  _T_945 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  _T_949 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  _T_953 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  _T_957 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  _T_961 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  _T_965 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  _T_969 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  _T_973 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  _T_977 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  _T_981 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  _T_985 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  _T_989 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  _T_993 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  _T_997 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  _T_1001 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  _T_1005 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  _T_1009 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  _T_1013 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  _T_1017 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  _T_1021 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  _T_1025 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  _T_1029 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  _T_1033 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  _T_1037 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  _T_1041 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  _T_1045 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  _T_1049 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  _T_1053 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  _T_1057 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  _T_1061 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  _T_1065 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  _T_1069 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  _T_1073 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  _T_1077 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  _T_1081 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  _T_1085 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  _T_1089 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  _T_1093 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  _T_1097 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  _T_1101 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  _T_1105 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  _T_1109 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  _T_1113 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  _T_1117 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  _T_1121 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  _T_1125 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  _T_1129 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  _T_1133 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  _T_1137 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  _T_1141 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  _T_1145 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  _T_1149 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  _T_1153 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  _T_1157 = _RAND_129[21:0];
  _RAND_130 = {1{`RANDOM}};
  _T_1161 = _RAND_130[21:0];
  _RAND_131 = {1{`RANDOM}};
  _T_1165 = _RAND_131[21:0];
  _RAND_132 = {1{`RANDOM}};
  _T_1169 = _RAND_132[21:0];
  _RAND_133 = {1{`RANDOM}};
  _T_1173 = _RAND_133[21:0];
  _RAND_134 = {1{`RANDOM}};
  _T_1177 = _RAND_134[21:0];
  _RAND_135 = {1{`RANDOM}};
  _T_1181 = _RAND_135[21:0];
  _RAND_136 = {1{`RANDOM}};
  _T_1185 = _RAND_136[21:0];
  _RAND_137 = {1{`RANDOM}};
  _T_1189 = _RAND_137[21:0];
  _RAND_138 = {1{`RANDOM}};
  _T_1193 = _RAND_138[21:0];
  _RAND_139 = {1{`RANDOM}};
  _T_1197 = _RAND_139[21:0];
  _RAND_140 = {1{`RANDOM}};
  _T_1201 = _RAND_140[21:0];
  _RAND_141 = {1{`RANDOM}};
  _T_1205 = _RAND_141[21:0];
  _RAND_142 = {1{`RANDOM}};
  _T_1209 = _RAND_142[21:0];
  _RAND_143 = {1{`RANDOM}};
  _T_1213 = _RAND_143[21:0];
  _RAND_144 = {1{`RANDOM}};
  _T_1217 = _RAND_144[21:0];
  _RAND_145 = {1{`RANDOM}};
  _T_1221 = _RAND_145[21:0];
  _RAND_146 = {1{`RANDOM}};
  _T_1225 = _RAND_146[21:0];
  _RAND_147 = {1{`RANDOM}};
  _T_1229 = _RAND_147[21:0];
  _RAND_148 = {1{`RANDOM}};
  _T_1233 = _RAND_148[21:0];
  _RAND_149 = {1{`RANDOM}};
  _T_1237 = _RAND_149[21:0];
  _RAND_150 = {1{`RANDOM}};
  _T_1241 = _RAND_150[21:0];
  _RAND_151 = {1{`RANDOM}};
  _T_1245 = _RAND_151[21:0];
  _RAND_152 = {1{`RANDOM}};
  _T_1249 = _RAND_152[21:0];
  _RAND_153 = {1{`RANDOM}};
  _T_1253 = _RAND_153[21:0];
  _RAND_154 = {1{`RANDOM}};
  _T_1257 = _RAND_154[21:0];
  _RAND_155 = {1{`RANDOM}};
  _T_1261 = _RAND_155[21:0];
  _RAND_156 = {1{`RANDOM}};
  _T_1265 = _RAND_156[21:0];
  _RAND_157 = {1{`RANDOM}};
  _T_1269 = _RAND_157[21:0];
  _RAND_158 = {1{`RANDOM}};
  _T_1273 = _RAND_158[21:0];
  _RAND_159 = {1{`RANDOM}};
  _T_1277 = _RAND_159[21:0];
  _RAND_160 = {1{`RANDOM}};
  _T_1281 = _RAND_160[21:0];
  _RAND_161 = {1{`RANDOM}};
  _T_1285 = _RAND_161[21:0];
  _RAND_162 = {1{`RANDOM}};
  _T_1289 = _RAND_162[21:0];
  _RAND_163 = {1{`RANDOM}};
  _T_1293 = _RAND_163[21:0];
  _RAND_164 = {1{`RANDOM}};
  _T_1297 = _RAND_164[21:0];
  _RAND_165 = {1{`RANDOM}};
  _T_1301 = _RAND_165[21:0];
  _RAND_166 = {1{`RANDOM}};
  _T_1305 = _RAND_166[21:0];
  _RAND_167 = {1{`RANDOM}};
  _T_1309 = _RAND_167[21:0];
  _RAND_168 = {1{`RANDOM}};
  _T_1313 = _RAND_168[21:0];
  _RAND_169 = {1{`RANDOM}};
  _T_1317 = _RAND_169[21:0];
  _RAND_170 = {1{`RANDOM}};
  _T_1321 = _RAND_170[21:0];
  _RAND_171 = {1{`RANDOM}};
  _T_1325 = _RAND_171[21:0];
  _RAND_172 = {1{`RANDOM}};
  _T_1329 = _RAND_172[21:0];
  _RAND_173 = {1{`RANDOM}};
  _T_1333 = _RAND_173[21:0];
  _RAND_174 = {1{`RANDOM}};
  _T_1337 = _RAND_174[21:0];
  _RAND_175 = {1{`RANDOM}};
  _T_1341 = _RAND_175[21:0];
  _RAND_176 = {1{`RANDOM}};
  _T_1345 = _RAND_176[21:0];
  _RAND_177 = {1{`RANDOM}};
  _T_1349 = _RAND_177[21:0];
  _RAND_178 = {1{`RANDOM}};
  _T_1353 = _RAND_178[21:0];
  _RAND_179 = {1{`RANDOM}};
  _T_1357 = _RAND_179[21:0];
  _RAND_180 = {1{`RANDOM}};
  _T_1361 = _RAND_180[21:0];
  _RAND_181 = {1{`RANDOM}};
  _T_1365 = _RAND_181[21:0];
  _RAND_182 = {1{`RANDOM}};
  _T_1369 = _RAND_182[21:0];
  _RAND_183 = {1{`RANDOM}};
  _T_1373 = _RAND_183[21:0];
  _RAND_184 = {1{`RANDOM}};
  _T_1377 = _RAND_184[21:0];
  _RAND_185 = {1{`RANDOM}};
  _T_1381 = _RAND_185[21:0];
  _RAND_186 = {1{`RANDOM}};
  _T_1385 = _RAND_186[21:0];
  _RAND_187 = {1{`RANDOM}};
  _T_1389 = _RAND_187[21:0];
  _RAND_188 = {1{`RANDOM}};
  _T_1393 = _RAND_188[21:0];
  _RAND_189 = {1{`RANDOM}};
  _T_1397 = _RAND_189[21:0];
  _RAND_190 = {1{`RANDOM}};
  _T_1401 = _RAND_190[21:0];
  _RAND_191 = {1{`RANDOM}};
  _T_1405 = _RAND_191[21:0];
  _RAND_192 = {1{`RANDOM}};
  _T_1409 = _RAND_192[21:0];
  _RAND_193 = {1{`RANDOM}};
  _T_1413 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  _T_1417 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  _T_1421 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  _T_1425 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  _T_1429 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  _T_1433 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  _T_1437 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  _T_1441 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  _T_1445 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  _T_1449 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  _T_1453 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  _T_1457 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  _T_1461 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  _T_1465 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  _T_1469 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  _T_1473 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  _T_1477 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  _T_1481 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  _T_1485 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  _T_1489 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  _T_1493 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  _T_1497 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  _T_1501 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  _T_1505 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  _T_1509 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  _T_1513 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  _T_1517 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  _T_1521 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  _T_1525 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  _T_1529 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  _T_1533 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  _T_1537 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  _T_1541 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  _T_1545 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  _T_1549 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  _T_1553 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  _T_1557 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  _T_1561 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  _T_1565 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  _T_1569 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  _T_1573 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  _T_1577 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  _T_1581 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  _T_1585 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  _T_1589 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  _T_1593 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  _T_1597 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  _T_1601 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  _T_1605 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  _T_1609 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  _T_1613 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  _T_1617 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  _T_1621 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  _T_1625 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  _T_1629 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  _T_1633 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  _T_1637 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  _T_1641 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  _T_1645 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  _T_1649 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  _T_1653 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  _T_1657 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  _T_1661 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  _T_1665 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  _T_1669 = _RAND_257[21:0];
  _RAND_258 = {1{`RANDOM}};
  _T_1673 = _RAND_258[21:0];
  _RAND_259 = {1{`RANDOM}};
  _T_1677 = _RAND_259[21:0];
  _RAND_260 = {1{`RANDOM}};
  _T_1681 = _RAND_260[21:0];
  _RAND_261 = {1{`RANDOM}};
  _T_1685 = _RAND_261[21:0];
  _RAND_262 = {1{`RANDOM}};
  _T_1689 = _RAND_262[21:0];
  _RAND_263 = {1{`RANDOM}};
  _T_1693 = _RAND_263[21:0];
  _RAND_264 = {1{`RANDOM}};
  _T_1697 = _RAND_264[21:0];
  _RAND_265 = {1{`RANDOM}};
  _T_1701 = _RAND_265[21:0];
  _RAND_266 = {1{`RANDOM}};
  _T_1705 = _RAND_266[21:0];
  _RAND_267 = {1{`RANDOM}};
  _T_1709 = _RAND_267[21:0];
  _RAND_268 = {1{`RANDOM}};
  _T_1713 = _RAND_268[21:0];
  _RAND_269 = {1{`RANDOM}};
  _T_1717 = _RAND_269[21:0];
  _RAND_270 = {1{`RANDOM}};
  _T_1721 = _RAND_270[21:0];
  _RAND_271 = {1{`RANDOM}};
  _T_1725 = _RAND_271[21:0];
  _RAND_272 = {1{`RANDOM}};
  _T_1729 = _RAND_272[21:0];
  _RAND_273 = {1{`RANDOM}};
  _T_1733 = _RAND_273[21:0];
  _RAND_274 = {1{`RANDOM}};
  _T_1737 = _RAND_274[21:0];
  _RAND_275 = {1{`RANDOM}};
  _T_1741 = _RAND_275[21:0];
  _RAND_276 = {1{`RANDOM}};
  _T_1745 = _RAND_276[21:0];
  _RAND_277 = {1{`RANDOM}};
  _T_1749 = _RAND_277[21:0];
  _RAND_278 = {1{`RANDOM}};
  _T_1753 = _RAND_278[21:0];
  _RAND_279 = {1{`RANDOM}};
  _T_1757 = _RAND_279[21:0];
  _RAND_280 = {1{`RANDOM}};
  _T_1761 = _RAND_280[21:0];
  _RAND_281 = {1{`RANDOM}};
  _T_1765 = _RAND_281[21:0];
  _RAND_282 = {1{`RANDOM}};
  _T_1769 = _RAND_282[21:0];
  _RAND_283 = {1{`RANDOM}};
  _T_1773 = _RAND_283[21:0];
  _RAND_284 = {1{`RANDOM}};
  _T_1777 = _RAND_284[21:0];
  _RAND_285 = {1{`RANDOM}};
  _T_1781 = _RAND_285[21:0];
  _RAND_286 = {1{`RANDOM}};
  _T_1785 = _RAND_286[21:0];
  _RAND_287 = {1{`RANDOM}};
  _T_1789 = _RAND_287[21:0];
  _RAND_288 = {1{`RANDOM}};
  _T_1793 = _RAND_288[21:0];
  _RAND_289 = {1{`RANDOM}};
  _T_1797 = _RAND_289[21:0];
  _RAND_290 = {1{`RANDOM}};
  _T_1801 = _RAND_290[21:0];
  _RAND_291 = {1{`RANDOM}};
  _T_1805 = _RAND_291[21:0];
  _RAND_292 = {1{`RANDOM}};
  _T_1809 = _RAND_292[21:0];
  _RAND_293 = {1{`RANDOM}};
  _T_1813 = _RAND_293[21:0];
  _RAND_294 = {1{`RANDOM}};
  _T_1817 = _RAND_294[21:0];
  _RAND_295 = {1{`RANDOM}};
  _T_1821 = _RAND_295[21:0];
  _RAND_296 = {1{`RANDOM}};
  _T_1825 = _RAND_296[21:0];
  _RAND_297 = {1{`RANDOM}};
  _T_1829 = _RAND_297[21:0];
  _RAND_298 = {1{`RANDOM}};
  _T_1833 = _RAND_298[21:0];
  _RAND_299 = {1{`RANDOM}};
  _T_1837 = _RAND_299[21:0];
  _RAND_300 = {1{`RANDOM}};
  _T_1841 = _RAND_300[21:0];
  _RAND_301 = {1{`RANDOM}};
  _T_1845 = _RAND_301[21:0];
  _RAND_302 = {1{`RANDOM}};
  _T_1849 = _RAND_302[21:0];
  _RAND_303 = {1{`RANDOM}};
  _T_1853 = _RAND_303[21:0];
  _RAND_304 = {1{`RANDOM}};
  _T_1857 = _RAND_304[21:0];
  _RAND_305 = {1{`RANDOM}};
  _T_1861 = _RAND_305[21:0];
  _RAND_306 = {1{`RANDOM}};
  _T_1865 = _RAND_306[21:0];
  _RAND_307 = {1{`RANDOM}};
  _T_1869 = _RAND_307[21:0];
  _RAND_308 = {1{`RANDOM}};
  _T_1873 = _RAND_308[21:0];
  _RAND_309 = {1{`RANDOM}};
  _T_1877 = _RAND_309[21:0];
  _RAND_310 = {1{`RANDOM}};
  _T_1881 = _RAND_310[21:0];
  _RAND_311 = {1{`RANDOM}};
  _T_1885 = _RAND_311[21:0];
  _RAND_312 = {1{`RANDOM}};
  _T_1889 = _RAND_312[21:0];
  _RAND_313 = {1{`RANDOM}};
  _T_1893 = _RAND_313[21:0];
  _RAND_314 = {1{`RANDOM}};
  _T_1897 = _RAND_314[21:0];
  _RAND_315 = {1{`RANDOM}};
  _T_1901 = _RAND_315[21:0];
  _RAND_316 = {1{`RANDOM}};
  _T_1905 = _RAND_316[21:0];
  _RAND_317 = {1{`RANDOM}};
  _T_1909 = _RAND_317[21:0];
  _RAND_318 = {1{`RANDOM}};
  _T_1913 = _RAND_318[21:0];
  _RAND_319 = {1{`RANDOM}};
  _T_1917 = _RAND_319[21:0];
  _RAND_320 = {1{`RANDOM}};
  _T_1921 = _RAND_320[21:0];
  _RAND_321 = {1{`RANDOM}};
  _T_1925 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  _T_1929 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  _T_1933 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  _T_1937 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  _T_1941 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  _T_1945 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  _T_1949 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  _T_1953 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  _T_1957 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  _T_1961 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  _T_1965 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  _T_1969 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  _T_1973 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  _T_1977 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  _T_1981 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  _T_1985 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  _T_1989 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  _T_1993 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  _T_1997 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  _T_2001 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  _T_2005 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  _T_2009 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  _T_2013 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  _T_2017 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  _T_2021 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  _T_2025 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  _T_2029 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  _T_2033 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  _T_2037 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  _T_2041 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  _T_2045 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  _T_2049 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  _T_2053 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  _T_2057 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  _T_2061 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  _T_2065 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  _T_2069 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  _T_2073 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  _T_2077 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  _T_2081 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  _T_2085 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  _T_2089 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  _T_2093 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  _T_2097 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  _T_2101 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  _T_2105 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  _T_2109 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  _T_2113 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  _T_2117 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  _T_2121 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  _T_2125 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  _T_2129 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  _T_2133 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  _T_2137 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  _T_2141 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  _T_2145 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  _T_2149 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  _T_2153 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  _T_2157 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  _T_2161 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  _T_2165 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  _T_2169 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  _T_2173 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  _T_2177 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  _T_2181 = _RAND_385[21:0];
  _RAND_386 = {1{`RANDOM}};
  _T_2185 = _RAND_386[21:0];
  _RAND_387 = {1{`RANDOM}};
  _T_2189 = _RAND_387[21:0];
  _RAND_388 = {1{`RANDOM}};
  _T_2193 = _RAND_388[21:0];
  _RAND_389 = {1{`RANDOM}};
  _T_2197 = _RAND_389[21:0];
  _RAND_390 = {1{`RANDOM}};
  _T_2201 = _RAND_390[21:0];
  _RAND_391 = {1{`RANDOM}};
  _T_2205 = _RAND_391[21:0];
  _RAND_392 = {1{`RANDOM}};
  _T_2209 = _RAND_392[21:0];
  _RAND_393 = {1{`RANDOM}};
  _T_2213 = _RAND_393[21:0];
  _RAND_394 = {1{`RANDOM}};
  _T_2217 = _RAND_394[21:0];
  _RAND_395 = {1{`RANDOM}};
  _T_2221 = _RAND_395[21:0];
  _RAND_396 = {1{`RANDOM}};
  _T_2225 = _RAND_396[21:0];
  _RAND_397 = {1{`RANDOM}};
  _T_2229 = _RAND_397[21:0];
  _RAND_398 = {1{`RANDOM}};
  _T_2233 = _RAND_398[21:0];
  _RAND_399 = {1{`RANDOM}};
  _T_2237 = _RAND_399[21:0];
  _RAND_400 = {1{`RANDOM}};
  _T_2241 = _RAND_400[21:0];
  _RAND_401 = {1{`RANDOM}};
  _T_2245 = _RAND_401[21:0];
  _RAND_402 = {1{`RANDOM}};
  _T_2249 = _RAND_402[21:0];
  _RAND_403 = {1{`RANDOM}};
  _T_2253 = _RAND_403[21:0];
  _RAND_404 = {1{`RANDOM}};
  _T_2257 = _RAND_404[21:0];
  _RAND_405 = {1{`RANDOM}};
  _T_2261 = _RAND_405[21:0];
  _RAND_406 = {1{`RANDOM}};
  _T_2265 = _RAND_406[21:0];
  _RAND_407 = {1{`RANDOM}};
  _T_2269 = _RAND_407[21:0];
  _RAND_408 = {1{`RANDOM}};
  _T_2273 = _RAND_408[21:0];
  _RAND_409 = {1{`RANDOM}};
  _T_2277 = _RAND_409[21:0];
  _RAND_410 = {1{`RANDOM}};
  _T_2281 = _RAND_410[21:0];
  _RAND_411 = {1{`RANDOM}};
  _T_2285 = _RAND_411[21:0];
  _RAND_412 = {1{`RANDOM}};
  _T_2289 = _RAND_412[21:0];
  _RAND_413 = {1{`RANDOM}};
  _T_2293 = _RAND_413[21:0];
  _RAND_414 = {1{`RANDOM}};
  _T_2297 = _RAND_414[21:0];
  _RAND_415 = {1{`RANDOM}};
  _T_2301 = _RAND_415[21:0];
  _RAND_416 = {1{`RANDOM}};
  _T_2305 = _RAND_416[21:0];
  _RAND_417 = {1{`RANDOM}};
  _T_2309 = _RAND_417[21:0];
  _RAND_418 = {1{`RANDOM}};
  _T_2313 = _RAND_418[21:0];
  _RAND_419 = {1{`RANDOM}};
  _T_2317 = _RAND_419[21:0];
  _RAND_420 = {1{`RANDOM}};
  _T_2321 = _RAND_420[21:0];
  _RAND_421 = {1{`RANDOM}};
  _T_2325 = _RAND_421[21:0];
  _RAND_422 = {1{`RANDOM}};
  _T_2329 = _RAND_422[21:0];
  _RAND_423 = {1{`RANDOM}};
  _T_2333 = _RAND_423[21:0];
  _RAND_424 = {1{`RANDOM}};
  _T_2337 = _RAND_424[21:0];
  _RAND_425 = {1{`RANDOM}};
  _T_2341 = _RAND_425[21:0];
  _RAND_426 = {1{`RANDOM}};
  _T_2345 = _RAND_426[21:0];
  _RAND_427 = {1{`RANDOM}};
  _T_2349 = _RAND_427[21:0];
  _RAND_428 = {1{`RANDOM}};
  _T_2353 = _RAND_428[21:0];
  _RAND_429 = {1{`RANDOM}};
  _T_2357 = _RAND_429[21:0];
  _RAND_430 = {1{`RANDOM}};
  _T_2361 = _RAND_430[21:0];
  _RAND_431 = {1{`RANDOM}};
  _T_2365 = _RAND_431[21:0];
  _RAND_432 = {1{`RANDOM}};
  _T_2369 = _RAND_432[21:0];
  _RAND_433 = {1{`RANDOM}};
  _T_2373 = _RAND_433[21:0];
  _RAND_434 = {1{`RANDOM}};
  _T_2377 = _RAND_434[21:0];
  _RAND_435 = {1{`RANDOM}};
  _T_2381 = _RAND_435[21:0];
  _RAND_436 = {1{`RANDOM}};
  _T_2385 = _RAND_436[21:0];
  _RAND_437 = {1{`RANDOM}};
  _T_2389 = _RAND_437[21:0];
  _RAND_438 = {1{`RANDOM}};
  _T_2393 = _RAND_438[21:0];
  _RAND_439 = {1{`RANDOM}};
  _T_2397 = _RAND_439[21:0];
  _RAND_440 = {1{`RANDOM}};
  _T_2401 = _RAND_440[21:0];
  _RAND_441 = {1{`RANDOM}};
  _T_2405 = _RAND_441[21:0];
  _RAND_442 = {1{`RANDOM}};
  _T_2409 = _RAND_442[21:0];
  _RAND_443 = {1{`RANDOM}};
  _T_2413 = _RAND_443[21:0];
  _RAND_444 = {1{`RANDOM}};
  _T_2417 = _RAND_444[21:0];
  _RAND_445 = {1{`RANDOM}};
  _T_2421 = _RAND_445[21:0];
  _RAND_446 = {1{`RANDOM}};
  _T_2425 = _RAND_446[21:0];
  _RAND_447 = {1{`RANDOM}};
  _T_2429 = _RAND_447[21:0];
  _RAND_448 = {1{`RANDOM}};
  _T_2433 = _RAND_448[21:0];
  _RAND_449 = {1{`RANDOM}};
  _T_2437 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  _T_2441 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  _T_2445 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  _T_2449 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  _T_2453 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  _T_2457 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  _T_2461 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  _T_2465 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  _T_2469 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  _T_2473 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  _T_2477 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  _T_2481 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  _T_2485 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  _T_2489 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  _T_2493 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  _T_2497 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  _T_2501 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  _T_2505 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  _T_2509 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  _T_2513 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  _T_2517 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  _T_2521 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  _T_2525 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  _T_2529 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  _T_2533 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  _T_2537 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  _T_2541 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  _T_2545 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  _T_2549 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  _T_2553 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  _T_2557 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  _T_2561 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  _T_2565 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  _T_2569 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  _T_2573 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  _T_2577 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  _T_2581 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  _T_2585 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  _T_2589 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  _T_2593 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  _T_2597 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  _T_2601 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  _T_2605 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  _T_2609 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  _T_2613 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  _T_2617 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  _T_2621 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  _T_2625 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  _T_2629 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  _T_2633 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  _T_2637 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  _T_2641 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  _T_2645 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  _T_2649 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  _T_2653 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  _T_2657 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  _T_2661 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  _T_2665 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  _T_2669 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  _T_2673 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  _T_2677 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  _T_2681 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  _T_2685 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  _T_2689 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  fghr = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_0 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_1 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_2 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_3 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_4 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_5 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_6 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_7 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_8 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_9 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_10 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_11 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_12 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_13 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_14 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_15 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_16 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_17 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_18 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_19 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_20 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_21 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_22 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_23 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_24 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_25 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_26 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_27 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_28 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_29 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_30 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_31 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_32 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_33 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_34 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_35 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_36 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_37 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_38 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_39 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_40 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_41 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_42 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_43 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_44 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_45 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_46 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_47 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_48 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_49 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_50 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_51 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_52 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_53 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_54 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_55 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_56 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_57 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_58 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_59 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_60 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_61 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_62 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_63 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_64 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_65 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_66 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_67 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_68 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_69 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_70 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_71 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_72 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_73 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_74 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_75 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_76 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_77 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_78 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_79 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_80 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_81 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_82 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_83 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_84 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_85 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_86 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_87 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_88 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_89 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_90 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_91 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_92 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_93 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_94 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_95 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_96 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_97 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_98 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_99 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_100 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_101 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_102 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_103 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_104 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_105 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_106 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_107 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_108 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_109 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_110 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_111 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_112 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_113 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_114 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_115 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_116 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_117 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_118 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_119 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_120 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_121 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_122 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_123 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_124 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_125 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_126 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_127 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_128 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_129 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_130 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_131 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_132 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_133 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_134 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_135 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_136 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_137 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_138 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_139 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_140 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_141 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_142 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_143 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_144 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_145 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_146 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_147 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_148 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_149 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_150 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_151 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_152 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_153 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_154 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_155 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_156 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_157 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_158 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_159 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_160 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_161 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_162 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_163 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_164 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_165 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_166 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_167 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_168 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_169 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_170 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_171 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_172 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_173 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_174 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_175 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_176 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_177 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_178 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_179 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_180 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_181 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_182 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_183 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_184 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_185 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_186 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_187 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_188 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_189 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_190 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_191 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_192 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_193 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_194 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_195 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_196 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_197 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_198 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_199 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_200 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_201 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_202 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_203 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_204 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_205 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_206 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_207 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_208 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_209 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_210 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_211 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_212 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_213 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_214 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_215 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_216 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_217 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_218 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_219 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_220 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_221 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_222 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_223 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_224 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_225 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_226 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_227 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_228 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_229 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_230 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_231 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_232 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_233 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_234 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_235 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_236 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_237 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_238 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_239 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_240 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_241 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_242 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_243 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_244 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_245 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_246 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_247 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_248 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_249 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_250 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_251 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_252 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_253 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_254 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_255 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_0 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_1 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_2 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_3 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_4 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_5 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_6 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_7 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_8 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_9 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_10 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_11 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_12 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_13 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_14 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_15 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_16 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_17 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_18 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_19 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_20 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_21 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_22 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_23 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_24 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_25 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_26 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_27 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_28 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_29 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_30 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_31 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_32 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_33 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_34 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_35 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_36 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_37 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_38 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_39 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_40 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_41 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_42 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_43 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_44 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_45 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_46 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_47 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_48 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_49 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_50 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_51 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_52 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_53 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_54 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_55 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_56 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_57 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_58 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_59 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_60 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_61 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_62 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_63 = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_64 = _RAND_834[1:0];
  _RAND_835 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_65 = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_66 = _RAND_836[1:0];
  _RAND_837 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_67 = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_68 = _RAND_838[1:0];
  _RAND_839 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_69 = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_70 = _RAND_840[1:0];
  _RAND_841 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_71 = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_72 = _RAND_842[1:0];
  _RAND_843 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_73 = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_74 = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_75 = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_76 = _RAND_846[1:0];
  _RAND_847 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_77 = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_78 = _RAND_848[1:0];
  _RAND_849 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_79 = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_80 = _RAND_850[1:0];
  _RAND_851 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_81 = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_82 = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_83 = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_84 = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_85 = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_86 = _RAND_856[1:0];
  _RAND_857 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_87 = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_88 = _RAND_858[1:0];
  _RAND_859 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_89 = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_90 = _RAND_860[1:0];
  _RAND_861 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_91 = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_92 = _RAND_862[1:0];
  _RAND_863 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_93 = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_94 = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_95 = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_96 = _RAND_866[1:0];
  _RAND_867 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_97 = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_98 = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_99 = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_100 = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_101 = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_102 = _RAND_872[1:0];
  _RAND_873 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_103 = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_104 = _RAND_874[1:0];
  _RAND_875 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_105 = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_106 = _RAND_876[1:0];
  _RAND_877 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_107 = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_108 = _RAND_878[1:0];
  _RAND_879 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_109 = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_110 = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_111 = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_112 = _RAND_882[1:0];
  _RAND_883 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_113 = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_114 = _RAND_884[1:0];
  _RAND_885 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_115 = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_116 = _RAND_886[1:0];
  _RAND_887 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_117 = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_118 = _RAND_888[1:0];
  _RAND_889 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_119 = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_120 = _RAND_890[1:0];
  _RAND_891 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_121 = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_122 = _RAND_892[1:0];
  _RAND_893 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_123 = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_124 = _RAND_894[1:0];
  _RAND_895 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_125 = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_126 = _RAND_896[1:0];
  _RAND_897 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_127 = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_128 = _RAND_898[1:0];
  _RAND_899 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_129 = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_130 = _RAND_900[1:0];
  _RAND_901 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_131 = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_132 = _RAND_902[1:0];
  _RAND_903 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_133 = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_134 = _RAND_904[1:0];
  _RAND_905 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_135 = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_136 = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_137 = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_138 = _RAND_908[1:0];
  _RAND_909 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_139 = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_140 = _RAND_910[1:0];
  _RAND_911 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_141 = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_142 = _RAND_912[1:0];
  _RAND_913 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_143 = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_144 = _RAND_914[1:0];
  _RAND_915 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_145 = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_146 = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_147 = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_148 = _RAND_918[1:0];
  _RAND_919 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_149 = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_150 = _RAND_920[1:0];
  _RAND_921 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_151 = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_152 = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_153 = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_154 = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_155 = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_156 = _RAND_926[1:0];
  _RAND_927 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_157 = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_158 = _RAND_928[1:0];
  _RAND_929 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_159 = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_160 = _RAND_930[1:0];
  _RAND_931 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_161 = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_162 = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_163 = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_164 = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_165 = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_166 = _RAND_936[1:0];
  _RAND_937 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_167 = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_168 = _RAND_938[1:0];
  _RAND_939 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_169 = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_170 = _RAND_940[1:0];
  _RAND_941 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_171 = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_172 = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_173 = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_174 = _RAND_944[1:0];
  _RAND_945 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_175 = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_176 = _RAND_946[1:0];
  _RAND_947 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_177 = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_178 = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_179 = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_180 = _RAND_950[1:0];
  _RAND_951 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_181 = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_182 = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_183 = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_184 = _RAND_954[1:0];
  _RAND_955 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_185 = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_186 = _RAND_956[1:0];
  _RAND_957 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_187 = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_188 = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_189 = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_190 = _RAND_960[1:0];
  _RAND_961 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_191 = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_192 = _RAND_962[1:0];
  _RAND_963 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_193 = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_194 = _RAND_964[1:0];
  _RAND_965 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_195 = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_196 = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_197 = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_198 = _RAND_968[1:0];
  _RAND_969 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_199 = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_200 = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_201 = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_202 = _RAND_972[1:0];
  _RAND_973 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_203 = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_204 = _RAND_974[1:0];
  _RAND_975 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_205 = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_206 = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_207 = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_208 = _RAND_978[1:0];
  _RAND_979 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_209 = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_210 = _RAND_980[1:0];
  _RAND_981 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_211 = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_212 = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_213 = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_214 = _RAND_984[1:0];
  _RAND_985 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_215 = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_216 = _RAND_986[1:0];
  _RAND_987 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_217 = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_218 = _RAND_988[1:0];
  _RAND_989 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_219 = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_220 = _RAND_990[1:0];
  _RAND_991 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_221 = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_222 = _RAND_992[1:0];
  _RAND_993 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_223 = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_224 = _RAND_994[1:0];
  _RAND_995 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_225 = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_226 = _RAND_996[1:0];
  _RAND_997 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_227 = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_228 = _RAND_998[1:0];
  _RAND_999 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_229 = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_230 = _RAND_1000[1:0];
  _RAND_1001 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_231 = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_232 = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_233 = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_234 = _RAND_1004[1:0];
  _RAND_1005 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_235 = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_236 = _RAND_1006[1:0];
  _RAND_1007 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_237 = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_238 = _RAND_1008[1:0];
  _RAND_1009 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_239 = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_240 = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_241 = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_242 = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_243 = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_244 = _RAND_1014[1:0];
  _RAND_1015 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_245 = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_246 = _RAND_1016[1:0];
  _RAND_1017 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_247 = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_248 = _RAND_1018[1:0];
  _RAND_1019 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_249 = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_250 = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_251 = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_252 = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_253 = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_254 = _RAND_1024[1:0];
  _RAND_1025 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_255 = _RAND_1025[1:0];
  _RAND_1026 = {1{`RANDOM}};
  exu_mp_way_f = _RAND_1026[0:0];
  _RAND_1027 = {8{`RANDOM}};
  btb_lru_b0_f = _RAND_1027[255:0];
  _RAND_1028 = {1{`RANDOM}};
  exu_flush_final_d1 = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  ifc_fetch_adder_prior = _RAND_1029[29:0];
  _RAND_1030 = {1{`RANDOM}};
  rets_out_0 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  rets_out_1 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  rets_out_2 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  rets_out_3 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  rets_out_4 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  rets_out_5 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  rets_out_6 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  rets_out_7 = _RAND_1037[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    leak_one_f_d1 = 1'h0;
  end
  if (reset) begin
    _T_645 = 22'h0;
  end
  if (reset) begin
    _T_649 = 22'h0;
  end
  if (reset) begin
    _T_653 = 22'h0;
  end
  if (reset) begin
    _T_657 = 22'h0;
  end
  if (reset) begin
    _T_661 = 22'h0;
  end
  if (reset) begin
    _T_665 = 22'h0;
  end
  if (reset) begin
    _T_669 = 22'h0;
  end
  if (reset) begin
    _T_673 = 22'h0;
  end
  if (reset) begin
    _T_677 = 22'h0;
  end
  if (reset) begin
    _T_681 = 22'h0;
  end
  if (reset) begin
    _T_685 = 22'h0;
  end
  if (reset) begin
    _T_689 = 22'h0;
  end
  if (reset) begin
    _T_693 = 22'h0;
  end
  if (reset) begin
    _T_697 = 22'h0;
  end
  if (reset) begin
    _T_701 = 22'h0;
  end
  if (reset) begin
    _T_705 = 22'h0;
  end
  if (reset) begin
    _T_709 = 22'h0;
  end
  if (reset) begin
    _T_713 = 22'h0;
  end
  if (reset) begin
    _T_717 = 22'h0;
  end
  if (reset) begin
    _T_721 = 22'h0;
  end
  if (reset) begin
    _T_725 = 22'h0;
  end
  if (reset) begin
    _T_729 = 22'h0;
  end
  if (reset) begin
    _T_733 = 22'h0;
  end
  if (reset) begin
    _T_737 = 22'h0;
  end
  if (reset) begin
    _T_741 = 22'h0;
  end
  if (reset) begin
    _T_745 = 22'h0;
  end
  if (reset) begin
    _T_749 = 22'h0;
  end
  if (reset) begin
    _T_753 = 22'h0;
  end
  if (reset) begin
    _T_757 = 22'h0;
  end
  if (reset) begin
    _T_761 = 22'h0;
  end
  if (reset) begin
    _T_765 = 22'h0;
  end
  if (reset) begin
    _T_769 = 22'h0;
  end
  if (reset) begin
    _T_773 = 22'h0;
  end
  if (reset) begin
    _T_777 = 22'h0;
  end
  if (reset) begin
    _T_781 = 22'h0;
  end
  if (reset) begin
    _T_785 = 22'h0;
  end
  if (reset) begin
    _T_789 = 22'h0;
  end
  if (reset) begin
    _T_793 = 22'h0;
  end
  if (reset) begin
    _T_797 = 22'h0;
  end
  if (reset) begin
    _T_801 = 22'h0;
  end
  if (reset) begin
    _T_805 = 22'h0;
  end
  if (reset) begin
    _T_809 = 22'h0;
  end
  if (reset) begin
    _T_813 = 22'h0;
  end
  if (reset) begin
    _T_817 = 22'h0;
  end
  if (reset) begin
    _T_821 = 22'h0;
  end
  if (reset) begin
    _T_825 = 22'h0;
  end
  if (reset) begin
    _T_829 = 22'h0;
  end
  if (reset) begin
    _T_833 = 22'h0;
  end
  if (reset) begin
    _T_837 = 22'h0;
  end
  if (reset) begin
    _T_841 = 22'h0;
  end
  if (reset) begin
    _T_845 = 22'h0;
  end
  if (reset) begin
    _T_849 = 22'h0;
  end
  if (reset) begin
    _T_853 = 22'h0;
  end
  if (reset) begin
    _T_857 = 22'h0;
  end
  if (reset) begin
    _T_861 = 22'h0;
  end
  if (reset) begin
    _T_865 = 22'h0;
  end
  if (reset) begin
    _T_869 = 22'h0;
  end
  if (reset) begin
    _T_873 = 22'h0;
  end
  if (reset) begin
    _T_877 = 22'h0;
  end
  if (reset) begin
    _T_881 = 22'h0;
  end
  if (reset) begin
    _T_885 = 22'h0;
  end
  if (reset) begin
    _T_889 = 22'h0;
  end
  if (reset) begin
    _T_893 = 22'h0;
  end
  if (reset) begin
    _T_897 = 22'h0;
  end
  if (reset) begin
    _T_901 = 22'h0;
  end
  if (reset) begin
    _T_905 = 22'h0;
  end
  if (reset) begin
    _T_909 = 22'h0;
  end
  if (reset) begin
    _T_913 = 22'h0;
  end
  if (reset) begin
    _T_917 = 22'h0;
  end
  if (reset) begin
    _T_921 = 22'h0;
  end
  if (reset) begin
    _T_925 = 22'h0;
  end
  if (reset) begin
    _T_929 = 22'h0;
  end
  if (reset) begin
    _T_933 = 22'h0;
  end
  if (reset) begin
    _T_937 = 22'h0;
  end
  if (reset) begin
    _T_941 = 22'h0;
  end
  if (reset) begin
    _T_945 = 22'h0;
  end
  if (reset) begin
    _T_949 = 22'h0;
  end
  if (reset) begin
    _T_953 = 22'h0;
  end
  if (reset) begin
    _T_957 = 22'h0;
  end
  if (reset) begin
    _T_961 = 22'h0;
  end
  if (reset) begin
    _T_965 = 22'h0;
  end
  if (reset) begin
    _T_969 = 22'h0;
  end
  if (reset) begin
    _T_973 = 22'h0;
  end
  if (reset) begin
    _T_977 = 22'h0;
  end
  if (reset) begin
    _T_981 = 22'h0;
  end
  if (reset) begin
    _T_985 = 22'h0;
  end
  if (reset) begin
    _T_989 = 22'h0;
  end
  if (reset) begin
    _T_993 = 22'h0;
  end
  if (reset) begin
    _T_997 = 22'h0;
  end
  if (reset) begin
    _T_1001 = 22'h0;
  end
  if (reset) begin
    _T_1005 = 22'h0;
  end
  if (reset) begin
    _T_1009 = 22'h0;
  end
  if (reset) begin
    _T_1013 = 22'h0;
  end
  if (reset) begin
    _T_1017 = 22'h0;
  end
  if (reset) begin
    _T_1021 = 22'h0;
  end
  if (reset) begin
    _T_1025 = 22'h0;
  end
  if (reset) begin
    _T_1029 = 22'h0;
  end
  if (reset) begin
    _T_1033 = 22'h0;
  end
  if (reset) begin
    _T_1037 = 22'h0;
  end
  if (reset) begin
    _T_1041 = 22'h0;
  end
  if (reset) begin
    _T_1045 = 22'h0;
  end
  if (reset) begin
    _T_1049 = 22'h0;
  end
  if (reset) begin
    _T_1053 = 22'h0;
  end
  if (reset) begin
    _T_1057 = 22'h0;
  end
  if (reset) begin
    _T_1061 = 22'h0;
  end
  if (reset) begin
    _T_1065 = 22'h0;
  end
  if (reset) begin
    _T_1069 = 22'h0;
  end
  if (reset) begin
    _T_1073 = 22'h0;
  end
  if (reset) begin
    _T_1077 = 22'h0;
  end
  if (reset) begin
    _T_1081 = 22'h0;
  end
  if (reset) begin
    _T_1085 = 22'h0;
  end
  if (reset) begin
    _T_1089 = 22'h0;
  end
  if (reset) begin
    _T_1093 = 22'h0;
  end
  if (reset) begin
    _T_1097 = 22'h0;
  end
  if (reset) begin
    _T_1101 = 22'h0;
  end
  if (reset) begin
    _T_1105 = 22'h0;
  end
  if (reset) begin
    _T_1109 = 22'h0;
  end
  if (reset) begin
    _T_1113 = 22'h0;
  end
  if (reset) begin
    _T_1117 = 22'h0;
  end
  if (reset) begin
    _T_1121 = 22'h0;
  end
  if (reset) begin
    _T_1125 = 22'h0;
  end
  if (reset) begin
    _T_1129 = 22'h0;
  end
  if (reset) begin
    _T_1133 = 22'h0;
  end
  if (reset) begin
    _T_1137 = 22'h0;
  end
  if (reset) begin
    _T_1141 = 22'h0;
  end
  if (reset) begin
    _T_1145 = 22'h0;
  end
  if (reset) begin
    _T_1149 = 22'h0;
  end
  if (reset) begin
    _T_1153 = 22'h0;
  end
  if (reset) begin
    _T_1157 = 22'h0;
  end
  if (reset) begin
    _T_1161 = 22'h0;
  end
  if (reset) begin
    _T_1165 = 22'h0;
  end
  if (reset) begin
    _T_1169 = 22'h0;
  end
  if (reset) begin
    _T_1173 = 22'h0;
  end
  if (reset) begin
    _T_1177 = 22'h0;
  end
  if (reset) begin
    _T_1181 = 22'h0;
  end
  if (reset) begin
    _T_1185 = 22'h0;
  end
  if (reset) begin
    _T_1189 = 22'h0;
  end
  if (reset) begin
    _T_1193 = 22'h0;
  end
  if (reset) begin
    _T_1197 = 22'h0;
  end
  if (reset) begin
    _T_1201 = 22'h0;
  end
  if (reset) begin
    _T_1205 = 22'h0;
  end
  if (reset) begin
    _T_1209 = 22'h0;
  end
  if (reset) begin
    _T_1213 = 22'h0;
  end
  if (reset) begin
    _T_1217 = 22'h0;
  end
  if (reset) begin
    _T_1221 = 22'h0;
  end
  if (reset) begin
    _T_1225 = 22'h0;
  end
  if (reset) begin
    _T_1229 = 22'h0;
  end
  if (reset) begin
    _T_1233 = 22'h0;
  end
  if (reset) begin
    _T_1237 = 22'h0;
  end
  if (reset) begin
    _T_1241 = 22'h0;
  end
  if (reset) begin
    _T_1245 = 22'h0;
  end
  if (reset) begin
    _T_1249 = 22'h0;
  end
  if (reset) begin
    _T_1253 = 22'h0;
  end
  if (reset) begin
    _T_1257 = 22'h0;
  end
  if (reset) begin
    _T_1261 = 22'h0;
  end
  if (reset) begin
    _T_1265 = 22'h0;
  end
  if (reset) begin
    _T_1269 = 22'h0;
  end
  if (reset) begin
    _T_1273 = 22'h0;
  end
  if (reset) begin
    _T_1277 = 22'h0;
  end
  if (reset) begin
    _T_1281 = 22'h0;
  end
  if (reset) begin
    _T_1285 = 22'h0;
  end
  if (reset) begin
    _T_1289 = 22'h0;
  end
  if (reset) begin
    _T_1293 = 22'h0;
  end
  if (reset) begin
    _T_1297 = 22'h0;
  end
  if (reset) begin
    _T_1301 = 22'h0;
  end
  if (reset) begin
    _T_1305 = 22'h0;
  end
  if (reset) begin
    _T_1309 = 22'h0;
  end
  if (reset) begin
    _T_1313 = 22'h0;
  end
  if (reset) begin
    _T_1317 = 22'h0;
  end
  if (reset) begin
    _T_1321 = 22'h0;
  end
  if (reset) begin
    _T_1325 = 22'h0;
  end
  if (reset) begin
    _T_1329 = 22'h0;
  end
  if (reset) begin
    _T_1333 = 22'h0;
  end
  if (reset) begin
    _T_1337 = 22'h0;
  end
  if (reset) begin
    _T_1341 = 22'h0;
  end
  if (reset) begin
    _T_1345 = 22'h0;
  end
  if (reset) begin
    _T_1349 = 22'h0;
  end
  if (reset) begin
    _T_1353 = 22'h0;
  end
  if (reset) begin
    _T_1357 = 22'h0;
  end
  if (reset) begin
    _T_1361 = 22'h0;
  end
  if (reset) begin
    _T_1365 = 22'h0;
  end
  if (reset) begin
    _T_1369 = 22'h0;
  end
  if (reset) begin
    _T_1373 = 22'h0;
  end
  if (reset) begin
    _T_1377 = 22'h0;
  end
  if (reset) begin
    _T_1381 = 22'h0;
  end
  if (reset) begin
    _T_1385 = 22'h0;
  end
  if (reset) begin
    _T_1389 = 22'h0;
  end
  if (reset) begin
    _T_1393 = 22'h0;
  end
  if (reset) begin
    _T_1397 = 22'h0;
  end
  if (reset) begin
    _T_1401 = 22'h0;
  end
  if (reset) begin
    _T_1405 = 22'h0;
  end
  if (reset) begin
    _T_1409 = 22'h0;
  end
  if (reset) begin
    _T_1413 = 22'h0;
  end
  if (reset) begin
    _T_1417 = 22'h0;
  end
  if (reset) begin
    _T_1421 = 22'h0;
  end
  if (reset) begin
    _T_1425 = 22'h0;
  end
  if (reset) begin
    _T_1429 = 22'h0;
  end
  if (reset) begin
    _T_1433 = 22'h0;
  end
  if (reset) begin
    _T_1437 = 22'h0;
  end
  if (reset) begin
    _T_1441 = 22'h0;
  end
  if (reset) begin
    _T_1445 = 22'h0;
  end
  if (reset) begin
    _T_1449 = 22'h0;
  end
  if (reset) begin
    _T_1453 = 22'h0;
  end
  if (reset) begin
    _T_1457 = 22'h0;
  end
  if (reset) begin
    _T_1461 = 22'h0;
  end
  if (reset) begin
    _T_1465 = 22'h0;
  end
  if (reset) begin
    _T_1469 = 22'h0;
  end
  if (reset) begin
    _T_1473 = 22'h0;
  end
  if (reset) begin
    _T_1477 = 22'h0;
  end
  if (reset) begin
    _T_1481 = 22'h0;
  end
  if (reset) begin
    _T_1485 = 22'h0;
  end
  if (reset) begin
    _T_1489 = 22'h0;
  end
  if (reset) begin
    _T_1493 = 22'h0;
  end
  if (reset) begin
    _T_1497 = 22'h0;
  end
  if (reset) begin
    _T_1501 = 22'h0;
  end
  if (reset) begin
    _T_1505 = 22'h0;
  end
  if (reset) begin
    _T_1509 = 22'h0;
  end
  if (reset) begin
    _T_1513 = 22'h0;
  end
  if (reset) begin
    _T_1517 = 22'h0;
  end
  if (reset) begin
    _T_1521 = 22'h0;
  end
  if (reset) begin
    _T_1525 = 22'h0;
  end
  if (reset) begin
    _T_1529 = 22'h0;
  end
  if (reset) begin
    _T_1533 = 22'h0;
  end
  if (reset) begin
    _T_1537 = 22'h0;
  end
  if (reset) begin
    _T_1541 = 22'h0;
  end
  if (reset) begin
    _T_1545 = 22'h0;
  end
  if (reset) begin
    _T_1549 = 22'h0;
  end
  if (reset) begin
    _T_1553 = 22'h0;
  end
  if (reset) begin
    _T_1557 = 22'h0;
  end
  if (reset) begin
    _T_1561 = 22'h0;
  end
  if (reset) begin
    _T_1565 = 22'h0;
  end
  if (reset) begin
    _T_1569 = 22'h0;
  end
  if (reset) begin
    _T_1573 = 22'h0;
  end
  if (reset) begin
    _T_1577 = 22'h0;
  end
  if (reset) begin
    _T_1581 = 22'h0;
  end
  if (reset) begin
    _T_1585 = 22'h0;
  end
  if (reset) begin
    _T_1589 = 22'h0;
  end
  if (reset) begin
    _T_1593 = 22'h0;
  end
  if (reset) begin
    _T_1597 = 22'h0;
  end
  if (reset) begin
    _T_1601 = 22'h0;
  end
  if (reset) begin
    _T_1605 = 22'h0;
  end
  if (reset) begin
    _T_1609 = 22'h0;
  end
  if (reset) begin
    _T_1613 = 22'h0;
  end
  if (reset) begin
    _T_1617 = 22'h0;
  end
  if (reset) begin
    _T_1621 = 22'h0;
  end
  if (reset) begin
    _T_1625 = 22'h0;
  end
  if (reset) begin
    _T_1629 = 22'h0;
  end
  if (reset) begin
    _T_1633 = 22'h0;
  end
  if (reset) begin
    _T_1637 = 22'h0;
  end
  if (reset) begin
    _T_1641 = 22'h0;
  end
  if (reset) begin
    _T_1645 = 22'h0;
  end
  if (reset) begin
    _T_1649 = 22'h0;
  end
  if (reset) begin
    _T_1653 = 22'h0;
  end
  if (reset) begin
    _T_1657 = 22'h0;
  end
  if (reset) begin
    _T_1661 = 22'h0;
  end
  if (reset) begin
    _T_1665 = 22'h0;
  end
  if (reset) begin
    _T_1669 = 22'h0;
  end
  if (reset) begin
    _T_1673 = 22'h0;
  end
  if (reset) begin
    _T_1677 = 22'h0;
  end
  if (reset) begin
    _T_1681 = 22'h0;
  end
  if (reset) begin
    _T_1685 = 22'h0;
  end
  if (reset) begin
    _T_1689 = 22'h0;
  end
  if (reset) begin
    _T_1693 = 22'h0;
  end
  if (reset) begin
    _T_1697 = 22'h0;
  end
  if (reset) begin
    _T_1701 = 22'h0;
  end
  if (reset) begin
    _T_1705 = 22'h0;
  end
  if (reset) begin
    _T_1709 = 22'h0;
  end
  if (reset) begin
    _T_1713 = 22'h0;
  end
  if (reset) begin
    _T_1717 = 22'h0;
  end
  if (reset) begin
    _T_1721 = 22'h0;
  end
  if (reset) begin
    _T_1725 = 22'h0;
  end
  if (reset) begin
    _T_1729 = 22'h0;
  end
  if (reset) begin
    _T_1733 = 22'h0;
  end
  if (reset) begin
    _T_1737 = 22'h0;
  end
  if (reset) begin
    _T_1741 = 22'h0;
  end
  if (reset) begin
    _T_1745 = 22'h0;
  end
  if (reset) begin
    _T_1749 = 22'h0;
  end
  if (reset) begin
    _T_1753 = 22'h0;
  end
  if (reset) begin
    _T_1757 = 22'h0;
  end
  if (reset) begin
    _T_1761 = 22'h0;
  end
  if (reset) begin
    _T_1765 = 22'h0;
  end
  if (reset) begin
    _T_1769 = 22'h0;
  end
  if (reset) begin
    _T_1773 = 22'h0;
  end
  if (reset) begin
    _T_1777 = 22'h0;
  end
  if (reset) begin
    _T_1781 = 22'h0;
  end
  if (reset) begin
    _T_1785 = 22'h0;
  end
  if (reset) begin
    _T_1789 = 22'h0;
  end
  if (reset) begin
    _T_1793 = 22'h0;
  end
  if (reset) begin
    _T_1797 = 22'h0;
  end
  if (reset) begin
    _T_1801 = 22'h0;
  end
  if (reset) begin
    _T_1805 = 22'h0;
  end
  if (reset) begin
    _T_1809 = 22'h0;
  end
  if (reset) begin
    _T_1813 = 22'h0;
  end
  if (reset) begin
    _T_1817 = 22'h0;
  end
  if (reset) begin
    _T_1821 = 22'h0;
  end
  if (reset) begin
    _T_1825 = 22'h0;
  end
  if (reset) begin
    _T_1829 = 22'h0;
  end
  if (reset) begin
    _T_1833 = 22'h0;
  end
  if (reset) begin
    _T_1837 = 22'h0;
  end
  if (reset) begin
    _T_1841 = 22'h0;
  end
  if (reset) begin
    _T_1845 = 22'h0;
  end
  if (reset) begin
    _T_1849 = 22'h0;
  end
  if (reset) begin
    _T_1853 = 22'h0;
  end
  if (reset) begin
    _T_1857 = 22'h0;
  end
  if (reset) begin
    _T_1861 = 22'h0;
  end
  if (reset) begin
    _T_1865 = 22'h0;
  end
  if (reset) begin
    _T_1869 = 22'h0;
  end
  if (reset) begin
    _T_1873 = 22'h0;
  end
  if (reset) begin
    _T_1877 = 22'h0;
  end
  if (reset) begin
    _T_1881 = 22'h0;
  end
  if (reset) begin
    _T_1885 = 22'h0;
  end
  if (reset) begin
    _T_1889 = 22'h0;
  end
  if (reset) begin
    _T_1893 = 22'h0;
  end
  if (reset) begin
    _T_1897 = 22'h0;
  end
  if (reset) begin
    _T_1901 = 22'h0;
  end
  if (reset) begin
    _T_1905 = 22'h0;
  end
  if (reset) begin
    _T_1909 = 22'h0;
  end
  if (reset) begin
    _T_1913 = 22'h0;
  end
  if (reset) begin
    _T_1917 = 22'h0;
  end
  if (reset) begin
    _T_1921 = 22'h0;
  end
  if (reset) begin
    _T_1925 = 22'h0;
  end
  if (reset) begin
    _T_1929 = 22'h0;
  end
  if (reset) begin
    _T_1933 = 22'h0;
  end
  if (reset) begin
    _T_1937 = 22'h0;
  end
  if (reset) begin
    _T_1941 = 22'h0;
  end
  if (reset) begin
    _T_1945 = 22'h0;
  end
  if (reset) begin
    _T_1949 = 22'h0;
  end
  if (reset) begin
    _T_1953 = 22'h0;
  end
  if (reset) begin
    _T_1957 = 22'h0;
  end
  if (reset) begin
    _T_1961 = 22'h0;
  end
  if (reset) begin
    _T_1965 = 22'h0;
  end
  if (reset) begin
    _T_1969 = 22'h0;
  end
  if (reset) begin
    _T_1973 = 22'h0;
  end
  if (reset) begin
    _T_1977 = 22'h0;
  end
  if (reset) begin
    _T_1981 = 22'h0;
  end
  if (reset) begin
    _T_1985 = 22'h0;
  end
  if (reset) begin
    _T_1989 = 22'h0;
  end
  if (reset) begin
    _T_1993 = 22'h0;
  end
  if (reset) begin
    _T_1997 = 22'h0;
  end
  if (reset) begin
    _T_2001 = 22'h0;
  end
  if (reset) begin
    _T_2005 = 22'h0;
  end
  if (reset) begin
    _T_2009 = 22'h0;
  end
  if (reset) begin
    _T_2013 = 22'h0;
  end
  if (reset) begin
    _T_2017 = 22'h0;
  end
  if (reset) begin
    _T_2021 = 22'h0;
  end
  if (reset) begin
    _T_2025 = 22'h0;
  end
  if (reset) begin
    _T_2029 = 22'h0;
  end
  if (reset) begin
    _T_2033 = 22'h0;
  end
  if (reset) begin
    _T_2037 = 22'h0;
  end
  if (reset) begin
    _T_2041 = 22'h0;
  end
  if (reset) begin
    _T_2045 = 22'h0;
  end
  if (reset) begin
    _T_2049 = 22'h0;
  end
  if (reset) begin
    _T_2053 = 22'h0;
  end
  if (reset) begin
    _T_2057 = 22'h0;
  end
  if (reset) begin
    _T_2061 = 22'h0;
  end
  if (reset) begin
    _T_2065 = 22'h0;
  end
  if (reset) begin
    _T_2069 = 22'h0;
  end
  if (reset) begin
    _T_2073 = 22'h0;
  end
  if (reset) begin
    _T_2077 = 22'h0;
  end
  if (reset) begin
    _T_2081 = 22'h0;
  end
  if (reset) begin
    _T_2085 = 22'h0;
  end
  if (reset) begin
    _T_2089 = 22'h0;
  end
  if (reset) begin
    _T_2093 = 22'h0;
  end
  if (reset) begin
    _T_2097 = 22'h0;
  end
  if (reset) begin
    _T_2101 = 22'h0;
  end
  if (reset) begin
    _T_2105 = 22'h0;
  end
  if (reset) begin
    _T_2109 = 22'h0;
  end
  if (reset) begin
    _T_2113 = 22'h0;
  end
  if (reset) begin
    _T_2117 = 22'h0;
  end
  if (reset) begin
    _T_2121 = 22'h0;
  end
  if (reset) begin
    _T_2125 = 22'h0;
  end
  if (reset) begin
    _T_2129 = 22'h0;
  end
  if (reset) begin
    _T_2133 = 22'h0;
  end
  if (reset) begin
    _T_2137 = 22'h0;
  end
  if (reset) begin
    _T_2141 = 22'h0;
  end
  if (reset) begin
    _T_2145 = 22'h0;
  end
  if (reset) begin
    _T_2149 = 22'h0;
  end
  if (reset) begin
    _T_2153 = 22'h0;
  end
  if (reset) begin
    _T_2157 = 22'h0;
  end
  if (reset) begin
    _T_2161 = 22'h0;
  end
  if (reset) begin
    _T_2165 = 22'h0;
  end
  if (reset) begin
    _T_2169 = 22'h0;
  end
  if (reset) begin
    _T_2173 = 22'h0;
  end
  if (reset) begin
    _T_2177 = 22'h0;
  end
  if (reset) begin
    _T_2181 = 22'h0;
  end
  if (reset) begin
    _T_2185 = 22'h0;
  end
  if (reset) begin
    _T_2189 = 22'h0;
  end
  if (reset) begin
    _T_2193 = 22'h0;
  end
  if (reset) begin
    _T_2197 = 22'h0;
  end
  if (reset) begin
    _T_2201 = 22'h0;
  end
  if (reset) begin
    _T_2205 = 22'h0;
  end
  if (reset) begin
    _T_2209 = 22'h0;
  end
  if (reset) begin
    _T_2213 = 22'h0;
  end
  if (reset) begin
    _T_2217 = 22'h0;
  end
  if (reset) begin
    _T_2221 = 22'h0;
  end
  if (reset) begin
    _T_2225 = 22'h0;
  end
  if (reset) begin
    _T_2229 = 22'h0;
  end
  if (reset) begin
    _T_2233 = 22'h0;
  end
  if (reset) begin
    _T_2237 = 22'h0;
  end
  if (reset) begin
    _T_2241 = 22'h0;
  end
  if (reset) begin
    _T_2245 = 22'h0;
  end
  if (reset) begin
    _T_2249 = 22'h0;
  end
  if (reset) begin
    _T_2253 = 22'h0;
  end
  if (reset) begin
    _T_2257 = 22'h0;
  end
  if (reset) begin
    _T_2261 = 22'h0;
  end
  if (reset) begin
    _T_2265 = 22'h0;
  end
  if (reset) begin
    _T_2269 = 22'h0;
  end
  if (reset) begin
    _T_2273 = 22'h0;
  end
  if (reset) begin
    _T_2277 = 22'h0;
  end
  if (reset) begin
    _T_2281 = 22'h0;
  end
  if (reset) begin
    _T_2285 = 22'h0;
  end
  if (reset) begin
    _T_2289 = 22'h0;
  end
  if (reset) begin
    _T_2293 = 22'h0;
  end
  if (reset) begin
    _T_2297 = 22'h0;
  end
  if (reset) begin
    _T_2301 = 22'h0;
  end
  if (reset) begin
    _T_2305 = 22'h0;
  end
  if (reset) begin
    _T_2309 = 22'h0;
  end
  if (reset) begin
    _T_2313 = 22'h0;
  end
  if (reset) begin
    _T_2317 = 22'h0;
  end
  if (reset) begin
    _T_2321 = 22'h0;
  end
  if (reset) begin
    _T_2325 = 22'h0;
  end
  if (reset) begin
    _T_2329 = 22'h0;
  end
  if (reset) begin
    _T_2333 = 22'h0;
  end
  if (reset) begin
    _T_2337 = 22'h0;
  end
  if (reset) begin
    _T_2341 = 22'h0;
  end
  if (reset) begin
    _T_2345 = 22'h0;
  end
  if (reset) begin
    _T_2349 = 22'h0;
  end
  if (reset) begin
    _T_2353 = 22'h0;
  end
  if (reset) begin
    _T_2357 = 22'h0;
  end
  if (reset) begin
    _T_2361 = 22'h0;
  end
  if (reset) begin
    _T_2365 = 22'h0;
  end
  if (reset) begin
    _T_2369 = 22'h0;
  end
  if (reset) begin
    _T_2373 = 22'h0;
  end
  if (reset) begin
    _T_2377 = 22'h0;
  end
  if (reset) begin
    _T_2381 = 22'h0;
  end
  if (reset) begin
    _T_2385 = 22'h0;
  end
  if (reset) begin
    _T_2389 = 22'h0;
  end
  if (reset) begin
    _T_2393 = 22'h0;
  end
  if (reset) begin
    _T_2397 = 22'h0;
  end
  if (reset) begin
    _T_2401 = 22'h0;
  end
  if (reset) begin
    _T_2405 = 22'h0;
  end
  if (reset) begin
    _T_2409 = 22'h0;
  end
  if (reset) begin
    _T_2413 = 22'h0;
  end
  if (reset) begin
    _T_2417 = 22'h0;
  end
  if (reset) begin
    _T_2421 = 22'h0;
  end
  if (reset) begin
    _T_2425 = 22'h0;
  end
  if (reset) begin
    _T_2429 = 22'h0;
  end
  if (reset) begin
    _T_2433 = 22'h0;
  end
  if (reset) begin
    _T_2437 = 22'h0;
  end
  if (reset) begin
    _T_2441 = 22'h0;
  end
  if (reset) begin
    _T_2445 = 22'h0;
  end
  if (reset) begin
    _T_2449 = 22'h0;
  end
  if (reset) begin
    _T_2453 = 22'h0;
  end
  if (reset) begin
    _T_2457 = 22'h0;
  end
  if (reset) begin
    _T_2461 = 22'h0;
  end
  if (reset) begin
    _T_2465 = 22'h0;
  end
  if (reset) begin
    _T_2469 = 22'h0;
  end
  if (reset) begin
    _T_2473 = 22'h0;
  end
  if (reset) begin
    _T_2477 = 22'h0;
  end
  if (reset) begin
    _T_2481 = 22'h0;
  end
  if (reset) begin
    _T_2485 = 22'h0;
  end
  if (reset) begin
    _T_2489 = 22'h0;
  end
  if (reset) begin
    _T_2493 = 22'h0;
  end
  if (reset) begin
    _T_2497 = 22'h0;
  end
  if (reset) begin
    _T_2501 = 22'h0;
  end
  if (reset) begin
    _T_2505 = 22'h0;
  end
  if (reset) begin
    _T_2509 = 22'h0;
  end
  if (reset) begin
    _T_2513 = 22'h0;
  end
  if (reset) begin
    _T_2517 = 22'h0;
  end
  if (reset) begin
    _T_2521 = 22'h0;
  end
  if (reset) begin
    _T_2525 = 22'h0;
  end
  if (reset) begin
    _T_2529 = 22'h0;
  end
  if (reset) begin
    _T_2533 = 22'h0;
  end
  if (reset) begin
    _T_2537 = 22'h0;
  end
  if (reset) begin
    _T_2541 = 22'h0;
  end
  if (reset) begin
    _T_2545 = 22'h0;
  end
  if (reset) begin
    _T_2549 = 22'h0;
  end
  if (reset) begin
    _T_2553 = 22'h0;
  end
  if (reset) begin
    _T_2557 = 22'h0;
  end
  if (reset) begin
    _T_2561 = 22'h0;
  end
  if (reset) begin
    _T_2565 = 22'h0;
  end
  if (reset) begin
    _T_2569 = 22'h0;
  end
  if (reset) begin
    _T_2573 = 22'h0;
  end
  if (reset) begin
    _T_2577 = 22'h0;
  end
  if (reset) begin
    _T_2581 = 22'h0;
  end
  if (reset) begin
    _T_2585 = 22'h0;
  end
  if (reset) begin
    _T_2589 = 22'h0;
  end
  if (reset) begin
    _T_2593 = 22'h0;
  end
  if (reset) begin
    _T_2597 = 22'h0;
  end
  if (reset) begin
    _T_2601 = 22'h0;
  end
  if (reset) begin
    _T_2605 = 22'h0;
  end
  if (reset) begin
    _T_2609 = 22'h0;
  end
  if (reset) begin
    _T_2613 = 22'h0;
  end
  if (reset) begin
    _T_2617 = 22'h0;
  end
  if (reset) begin
    _T_2621 = 22'h0;
  end
  if (reset) begin
    _T_2625 = 22'h0;
  end
  if (reset) begin
    _T_2629 = 22'h0;
  end
  if (reset) begin
    _T_2633 = 22'h0;
  end
  if (reset) begin
    _T_2637 = 22'h0;
  end
  if (reset) begin
    _T_2641 = 22'h0;
  end
  if (reset) begin
    _T_2645 = 22'h0;
  end
  if (reset) begin
    _T_2649 = 22'h0;
  end
  if (reset) begin
    _T_2653 = 22'h0;
  end
  if (reset) begin
    _T_2657 = 22'h0;
  end
  if (reset) begin
    _T_2661 = 22'h0;
  end
  if (reset) begin
    _T_2665 = 22'h0;
  end
  if (reset) begin
    _T_2669 = 22'h0;
  end
  if (reset) begin
    _T_2673 = 22'h0;
  end
  if (reset) begin
    _T_2677 = 22'h0;
  end
  if (reset) begin
    _T_2681 = 22'h0;
  end
  if (reset) begin
    _T_2685 = 22'h0;
  end
  if (reset) begin
    _T_2689 = 22'h0;
  end
  if (reset) begin
    fghr = 8'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_255 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_255 = 2'h0;
  end
  if (reset) begin
    exu_mp_way_f = 1'h0;
  end
  if (reset) begin
    btb_lru_b0_f = 256'h0;
  end
  if (reset) begin
    exu_flush_final_d1 = 1'h0;
  end
  if (reset) begin
    ifc_fetch_adder_prior = 30'h0;
  end
  if (reset) begin
    rets_out_0 = 32'h0;
  end
  if (reset) begin
    rets_out_1 = 32'h0;
  end
  if (reset) begin
    rets_out_2 = 32'h0;
  end
  if (reset) begin
    rets_out_3 = 32'h0;
  end
  if (reset) begin
    rets_out_4 = 32'h0;
  end
  if (reset) begin
    rets_out_5 = 32'h0;
  end
  if (reset) begin
    rets_out_6 = 32'h0;
  end
  if (reset) begin
    rets_out_7 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      leak_one_f_d1 <= 1'h0;
    end else if (_T_363) begin
      leak_one_f_d1 <= leak_one_f;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_645 <= 22'h0;
    end else if (_T_643) begin
      _T_645 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_649 <= 22'h0;
    end else if (_T_647) begin
      _T_649 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_653 <= 22'h0;
    end else if (_T_651) begin
      _T_653 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_657 <= 22'h0;
    end else if (_T_655) begin
      _T_657 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_661 <= 22'h0;
    end else if (_T_659) begin
      _T_661 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_665 <= 22'h0;
    end else if (_T_663) begin
      _T_665 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_669 <= 22'h0;
    end else if (_T_667) begin
      _T_669 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_673 <= 22'h0;
    end else if (_T_671) begin
      _T_673 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_677 <= 22'h0;
    end else if (_T_675) begin
      _T_677 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_681 <= 22'h0;
    end else if (_T_679) begin
      _T_681 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_685 <= 22'h0;
    end else if (_T_683) begin
      _T_685 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_689 <= 22'h0;
    end else if (_T_687) begin
      _T_689 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_693 <= 22'h0;
    end else if (_T_691) begin
      _T_693 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_697 <= 22'h0;
    end else if (_T_695) begin
      _T_697 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_701 <= 22'h0;
    end else if (_T_699) begin
      _T_701 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_705 <= 22'h0;
    end else if (_T_703) begin
      _T_705 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_709 <= 22'h0;
    end else if (_T_707) begin
      _T_709 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_713 <= 22'h0;
    end else if (_T_711) begin
      _T_713 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_717 <= 22'h0;
    end else if (_T_715) begin
      _T_717 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_721 <= 22'h0;
    end else if (_T_719) begin
      _T_721 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_725 <= 22'h0;
    end else if (_T_723) begin
      _T_725 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_729 <= 22'h0;
    end else if (_T_727) begin
      _T_729 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_733 <= 22'h0;
    end else if (_T_731) begin
      _T_733 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_737 <= 22'h0;
    end else if (_T_735) begin
      _T_737 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_741 <= 22'h0;
    end else if (_T_739) begin
      _T_741 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_745 <= 22'h0;
    end else if (_T_743) begin
      _T_745 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_749 <= 22'h0;
    end else if (_T_747) begin
      _T_749 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_753 <= 22'h0;
    end else if (_T_751) begin
      _T_753 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_757 <= 22'h0;
    end else if (_T_755) begin
      _T_757 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_761 <= 22'h0;
    end else if (_T_759) begin
      _T_761 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_765 <= 22'h0;
    end else if (_T_763) begin
      _T_765 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_769 <= 22'h0;
    end else if (_T_767) begin
      _T_769 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_773 <= 22'h0;
    end else if (_T_771) begin
      _T_773 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_777 <= 22'h0;
    end else if (_T_775) begin
      _T_777 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_781 <= 22'h0;
    end else if (_T_779) begin
      _T_781 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_785 <= 22'h0;
    end else if (_T_783) begin
      _T_785 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_789 <= 22'h0;
    end else if (_T_787) begin
      _T_789 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_793 <= 22'h0;
    end else if (_T_791) begin
      _T_793 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_797 <= 22'h0;
    end else if (_T_795) begin
      _T_797 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_801 <= 22'h0;
    end else if (_T_799) begin
      _T_801 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_805 <= 22'h0;
    end else if (_T_803) begin
      _T_805 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_809 <= 22'h0;
    end else if (_T_807) begin
      _T_809 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_813 <= 22'h0;
    end else if (_T_811) begin
      _T_813 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_817 <= 22'h0;
    end else if (_T_815) begin
      _T_817 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_821 <= 22'h0;
    end else if (_T_819) begin
      _T_821 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_825 <= 22'h0;
    end else if (_T_823) begin
      _T_825 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_829 <= 22'h0;
    end else if (_T_827) begin
      _T_829 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_833 <= 22'h0;
    end else if (_T_831) begin
      _T_833 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_837 <= 22'h0;
    end else if (_T_835) begin
      _T_837 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_841 <= 22'h0;
    end else if (_T_839) begin
      _T_841 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_845 <= 22'h0;
    end else if (_T_843) begin
      _T_845 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_849 <= 22'h0;
    end else if (_T_847) begin
      _T_849 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_853 <= 22'h0;
    end else if (_T_851) begin
      _T_853 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_857 <= 22'h0;
    end else if (_T_855) begin
      _T_857 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_861 <= 22'h0;
    end else if (_T_859) begin
      _T_861 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_865 <= 22'h0;
    end else if (_T_863) begin
      _T_865 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_869 <= 22'h0;
    end else if (_T_867) begin
      _T_869 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_873 <= 22'h0;
    end else if (_T_871) begin
      _T_873 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_877 <= 22'h0;
    end else if (_T_875) begin
      _T_877 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_881 <= 22'h0;
    end else if (_T_879) begin
      _T_881 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_885 <= 22'h0;
    end else if (_T_883) begin
      _T_885 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_889 <= 22'h0;
    end else if (_T_887) begin
      _T_889 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_893 <= 22'h0;
    end else if (_T_891) begin
      _T_893 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_897 <= 22'h0;
    end else if (_T_895) begin
      _T_897 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_901 <= 22'h0;
    end else if (_T_899) begin
      _T_901 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_905 <= 22'h0;
    end else if (_T_903) begin
      _T_905 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_909 <= 22'h0;
    end else if (_T_907) begin
      _T_909 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_913 <= 22'h0;
    end else if (_T_911) begin
      _T_913 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_917 <= 22'h0;
    end else if (_T_915) begin
      _T_917 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_921 <= 22'h0;
    end else if (_T_919) begin
      _T_921 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_925 <= 22'h0;
    end else if (_T_923) begin
      _T_925 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_929 <= 22'h0;
    end else if (_T_927) begin
      _T_929 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_933 <= 22'h0;
    end else if (_T_931) begin
      _T_933 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_937 <= 22'h0;
    end else if (_T_935) begin
      _T_937 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_941 <= 22'h0;
    end else if (_T_939) begin
      _T_941 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_945 <= 22'h0;
    end else if (_T_943) begin
      _T_945 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_949 <= 22'h0;
    end else if (_T_947) begin
      _T_949 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_953 <= 22'h0;
    end else if (_T_951) begin
      _T_953 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_957 <= 22'h0;
    end else if (_T_955) begin
      _T_957 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_961 <= 22'h0;
    end else if (_T_959) begin
      _T_961 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_965 <= 22'h0;
    end else if (_T_963) begin
      _T_965 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_969 <= 22'h0;
    end else if (_T_967) begin
      _T_969 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_973 <= 22'h0;
    end else if (_T_971) begin
      _T_973 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_977 <= 22'h0;
    end else if (_T_975) begin
      _T_977 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_981 <= 22'h0;
    end else if (_T_979) begin
      _T_981 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_985 <= 22'h0;
    end else if (_T_983) begin
      _T_985 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_989 <= 22'h0;
    end else if (_T_987) begin
      _T_989 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_993 <= 22'h0;
    end else if (_T_991) begin
      _T_993 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_997 <= 22'h0;
    end else if (_T_995) begin
      _T_997 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1001 <= 22'h0;
    end else if (_T_999) begin
      _T_1001 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1005 <= 22'h0;
    end else if (_T_1003) begin
      _T_1005 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1009 <= 22'h0;
    end else if (_T_1007) begin
      _T_1009 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1013 <= 22'h0;
    end else if (_T_1011) begin
      _T_1013 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1017 <= 22'h0;
    end else if (_T_1015) begin
      _T_1017 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1021 <= 22'h0;
    end else if (_T_1019) begin
      _T_1021 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1025 <= 22'h0;
    end else if (_T_1023) begin
      _T_1025 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1029 <= 22'h0;
    end else if (_T_1027) begin
      _T_1029 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1033 <= 22'h0;
    end else if (_T_1031) begin
      _T_1033 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1037 <= 22'h0;
    end else if (_T_1035) begin
      _T_1037 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1041 <= 22'h0;
    end else if (_T_1039) begin
      _T_1041 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1045 <= 22'h0;
    end else if (_T_1043) begin
      _T_1045 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1049 <= 22'h0;
    end else if (_T_1047) begin
      _T_1049 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1053 <= 22'h0;
    end else if (_T_1051) begin
      _T_1053 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1057 <= 22'h0;
    end else if (_T_1055) begin
      _T_1057 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1061 <= 22'h0;
    end else if (_T_1059) begin
      _T_1061 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1065 <= 22'h0;
    end else if (_T_1063) begin
      _T_1065 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1069 <= 22'h0;
    end else if (_T_1067) begin
      _T_1069 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1073 <= 22'h0;
    end else if (_T_1071) begin
      _T_1073 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1077 <= 22'h0;
    end else if (_T_1075) begin
      _T_1077 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1081 <= 22'h0;
    end else if (_T_1079) begin
      _T_1081 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1085 <= 22'h0;
    end else if (_T_1083) begin
      _T_1085 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1089 <= 22'h0;
    end else if (_T_1087) begin
      _T_1089 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1093 <= 22'h0;
    end else if (_T_1091) begin
      _T_1093 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1097 <= 22'h0;
    end else if (_T_1095) begin
      _T_1097 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1101 <= 22'h0;
    end else if (_T_1099) begin
      _T_1101 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1105 <= 22'h0;
    end else if (_T_1103) begin
      _T_1105 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1109 <= 22'h0;
    end else if (_T_1107) begin
      _T_1109 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1113 <= 22'h0;
    end else if (_T_1111) begin
      _T_1113 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1117 <= 22'h0;
    end else if (_T_1115) begin
      _T_1117 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1121 <= 22'h0;
    end else if (_T_1119) begin
      _T_1121 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1125 <= 22'h0;
    end else if (_T_1123) begin
      _T_1125 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1129 <= 22'h0;
    end else if (_T_1127) begin
      _T_1129 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1133 <= 22'h0;
    end else if (_T_1131) begin
      _T_1133 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1137 <= 22'h0;
    end else if (_T_1135) begin
      _T_1137 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1141 <= 22'h0;
    end else if (_T_1139) begin
      _T_1141 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1145 <= 22'h0;
    end else if (_T_1143) begin
      _T_1145 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1149 <= 22'h0;
    end else if (_T_1147) begin
      _T_1149 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1153 <= 22'h0;
    end else if (_T_1151) begin
      _T_1153 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1157 <= 22'h0;
    end else if (_T_1155) begin
      _T_1157 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1161 <= 22'h0;
    end else if (_T_1159) begin
      _T_1161 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1165 <= 22'h0;
    end else if (_T_1163) begin
      _T_1165 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1169 <= 22'h0;
    end else if (_T_1167) begin
      _T_1169 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1173 <= 22'h0;
    end else if (_T_1171) begin
      _T_1173 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1177 <= 22'h0;
    end else if (_T_1175) begin
      _T_1177 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1181 <= 22'h0;
    end else if (_T_1179) begin
      _T_1181 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1185 <= 22'h0;
    end else if (_T_1183) begin
      _T_1185 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1189 <= 22'h0;
    end else if (_T_1187) begin
      _T_1189 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1193 <= 22'h0;
    end else if (_T_1191) begin
      _T_1193 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1197 <= 22'h0;
    end else if (_T_1195) begin
      _T_1197 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1201 <= 22'h0;
    end else if (_T_1199) begin
      _T_1201 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1205 <= 22'h0;
    end else if (_T_1203) begin
      _T_1205 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1209 <= 22'h0;
    end else if (_T_1207) begin
      _T_1209 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1213 <= 22'h0;
    end else if (_T_1211) begin
      _T_1213 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1217 <= 22'h0;
    end else if (_T_1215) begin
      _T_1217 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1221 <= 22'h0;
    end else if (_T_1219) begin
      _T_1221 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1225 <= 22'h0;
    end else if (_T_1223) begin
      _T_1225 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1229 <= 22'h0;
    end else if (_T_1227) begin
      _T_1229 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1233 <= 22'h0;
    end else if (_T_1231) begin
      _T_1233 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1237 <= 22'h0;
    end else if (_T_1235) begin
      _T_1237 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1241 <= 22'h0;
    end else if (_T_1239) begin
      _T_1241 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1245 <= 22'h0;
    end else if (_T_1243) begin
      _T_1245 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1249 <= 22'h0;
    end else if (_T_1247) begin
      _T_1249 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1253 <= 22'h0;
    end else if (_T_1251) begin
      _T_1253 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1257 <= 22'h0;
    end else if (_T_1255) begin
      _T_1257 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1261 <= 22'h0;
    end else if (_T_1259) begin
      _T_1261 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1265 <= 22'h0;
    end else if (_T_1263) begin
      _T_1265 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1269 <= 22'h0;
    end else if (_T_1267) begin
      _T_1269 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1273 <= 22'h0;
    end else if (_T_1271) begin
      _T_1273 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1277 <= 22'h0;
    end else if (_T_1275) begin
      _T_1277 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1281 <= 22'h0;
    end else if (_T_1279) begin
      _T_1281 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1285 <= 22'h0;
    end else if (_T_1283) begin
      _T_1285 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1289 <= 22'h0;
    end else if (_T_1287) begin
      _T_1289 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1293 <= 22'h0;
    end else if (_T_1291) begin
      _T_1293 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1297 <= 22'h0;
    end else if (_T_1295) begin
      _T_1297 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1301 <= 22'h0;
    end else if (_T_1299) begin
      _T_1301 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1305 <= 22'h0;
    end else if (_T_1303) begin
      _T_1305 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1309 <= 22'h0;
    end else if (_T_1307) begin
      _T_1309 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1313 <= 22'h0;
    end else if (_T_1311) begin
      _T_1313 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1317 <= 22'h0;
    end else if (_T_1315) begin
      _T_1317 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1321 <= 22'h0;
    end else if (_T_1319) begin
      _T_1321 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1325 <= 22'h0;
    end else if (_T_1323) begin
      _T_1325 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1329 <= 22'h0;
    end else if (_T_1327) begin
      _T_1329 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1333 <= 22'h0;
    end else if (_T_1331) begin
      _T_1333 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1337 <= 22'h0;
    end else if (_T_1335) begin
      _T_1337 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1341 <= 22'h0;
    end else if (_T_1339) begin
      _T_1341 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1345 <= 22'h0;
    end else if (_T_1343) begin
      _T_1345 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1349 <= 22'h0;
    end else if (_T_1347) begin
      _T_1349 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1353 <= 22'h0;
    end else if (_T_1351) begin
      _T_1353 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1357 <= 22'h0;
    end else if (_T_1355) begin
      _T_1357 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1361 <= 22'h0;
    end else if (_T_1359) begin
      _T_1361 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1365 <= 22'h0;
    end else if (_T_1363) begin
      _T_1365 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1369 <= 22'h0;
    end else if (_T_1367) begin
      _T_1369 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1373 <= 22'h0;
    end else if (_T_1371) begin
      _T_1373 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1377 <= 22'h0;
    end else if (_T_1375) begin
      _T_1377 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1381 <= 22'h0;
    end else if (_T_1379) begin
      _T_1381 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1385 <= 22'h0;
    end else if (_T_1383) begin
      _T_1385 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1389 <= 22'h0;
    end else if (_T_1387) begin
      _T_1389 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1393 <= 22'h0;
    end else if (_T_1391) begin
      _T_1393 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1397 <= 22'h0;
    end else if (_T_1395) begin
      _T_1397 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1401 <= 22'h0;
    end else if (_T_1399) begin
      _T_1401 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1405 <= 22'h0;
    end else if (_T_1403) begin
      _T_1405 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1409 <= 22'h0;
    end else if (_T_1407) begin
      _T_1409 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1413 <= 22'h0;
    end else if (_T_1411) begin
      _T_1413 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1417 <= 22'h0;
    end else if (_T_1415) begin
      _T_1417 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1421 <= 22'h0;
    end else if (_T_1419) begin
      _T_1421 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1425 <= 22'h0;
    end else if (_T_1423) begin
      _T_1425 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1429 <= 22'h0;
    end else if (_T_1427) begin
      _T_1429 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1433 <= 22'h0;
    end else if (_T_1431) begin
      _T_1433 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1437 <= 22'h0;
    end else if (_T_1435) begin
      _T_1437 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1441 <= 22'h0;
    end else if (_T_1439) begin
      _T_1441 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1445 <= 22'h0;
    end else if (_T_1443) begin
      _T_1445 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1449 <= 22'h0;
    end else if (_T_1447) begin
      _T_1449 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1453 <= 22'h0;
    end else if (_T_1451) begin
      _T_1453 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1457 <= 22'h0;
    end else if (_T_1455) begin
      _T_1457 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1461 <= 22'h0;
    end else if (_T_1459) begin
      _T_1461 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1465 <= 22'h0;
    end else if (_T_1463) begin
      _T_1465 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1469 <= 22'h0;
    end else if (_T_1467) begin
      _T_1469 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1473 <= 22'h0;
    end else if (_T_1471) begin
      _T_1473 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1477 <= 22'h0;
    end else if (_T_1475) begin
      _T_1477 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1481 <= 22'h0;
    end else if (_T_1479) begin
      _T_1481 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1485 <= 22'h0;
    end else if (_T_1483) begin
      _T_1485 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1489 <= 22'h0;
    end else if (_T_1487) begin
      _T_1489 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1493 <= 22'h0;
    end else if (_T_1491) begin
      _T_1493 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1497 <= 22'h0;
    end else if (_T_1495) begin
      _T_1497 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1501 <= 22'h0;
    end else if (_T_1499) begin
      _T_1501 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1505 <= 22'h0;
    end else if (_T_1503) begin
      _T_1505 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1509 <= 22'h0;
    end else if (_T_1507) begin
      _T_1509 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1513 <= 22'h0;
    end else if (_T_1511) begin
      _T_1513 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1517 <= 22'h0;
    end else if (_T_1515) begin
      _T_1517 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1521 <= 22'h0;
    end else if (_T_1519) begin
      _T_1521 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1525 <= 22'h0;
    end else if (_T_1523) begin
      _T_1525 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1529 <= 22'h0;
    end else if (_T_1527) begin
      _T_1529 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1533 <= 22'h0;
    end else if (_T_1531) begin
      _T_1533 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1537 <= 22'h0;
    end else if (_T_1535) begin
      _T_1537 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1541 <= 22'h0;
    end else if (_T_1539) begin
      _T_1541 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1545 <= 22'h0;
    end else if (_T_1543) begin
      _T_1545 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1549 <= 22'h0;
    end else if (_T_1547) begin
      _T_1549 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1553 <= 22'h0;
    end else if (_T_1551) begin
      _T_1553 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1557 <= 22'h0;
    end else if (_T_1555) begin
      _T_1557 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1561 <= 22'h0;
    end else if (_T_1559) begin
      _T_1561 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1565 <= 22'h0;
    end else if (_T_1563) begin
      _T_1565 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1569 <= 22'h0;
    end else if (_T_1567) begin
      _T_1569 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1573 <= 22'h0;
    end else if (_T_1571) begin
      _T_1573 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1577 <= 22'h0;
    end else if (_T_1575) begin
      _T_1577 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1581 <= 22'h0;
    end else if (_T_1579) begin
      _T_1581 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1585 <= 22'h0;
    end else if (_T_1583) begin
      _T_1585 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1589 <= 22'h0;
    end else if (_T_1587) begin
      _T_1589 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1593 <= 22'h0;
    end else if (_T_1591) begin
      _T_1593 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1597 <= 22'h0;
    end else if (_T_1595) begin
      _T_1597 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1601 <= 22'h0;
    end else if (_T_1599) begin
      _T_1601 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1605 <= 22'h0;
    end else if (_T_1603) begin
      _T_1605 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1609 <= 22'h0;
    end else if (_T_1607) begin
      _T_1609 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1613 <= 22'h0;
    end else if (_T_1611) begin
      _T_1613 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1617 <= 22'h0;
    end else if (_T_1615) begin
      _T_1617 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1621 <= 22'h0;
    end else if (_T_1619) begin
      _T_1621 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1625 <= 22'h0;
    end else if (_T_1623) begin
      _T_1625 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1629 <= 22'h0;
    end else if (_T_1627) begin
      _T_1629 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1633 <= 22'h0;
    end else if (_T_1631) begin
      _T_1633 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1637 <= 22'h0;
    end else if (_T_1635) begin
      _T_1637 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1641 <= 22'h0;
    end else if (_T_1639) begin
      _T_1641 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1645 <= 22'h0;
    end else if (_T_1643) begin
      _T_1645 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1649 <= 22'h0;
    end else if (_T_1647) begin
      _T_1649 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1653 <= 22'h0;
    end else if (_T_1651) begin
      _T_1653 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1657 <= 22'h0;
    end else if (_T_1655) begin
      _T_1657 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1661 <= 22'h0;
    end else if (_T_1659) begin
      _T_1661 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1665 <= 22'h0;
    end else if (_T_1663) begin
      _T_1665 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1669 <= 22'h0;
    end else if (_T_1667) begin
      _T_1669 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1673 <= 22'h0;
    end else if (_T_1671) begin
      _T_1673 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1677 <= 22'h0;
    end else if (_T_1675) begin
      _T_1677 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1681 <= 22'h0;
    end else if (_T_1679) begin
      _T_1681 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1685 <= 22'h0;
    end else if (_T_1683) begin
      _T_1685 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1689 <= 22'h0;
    end else if (_T_1687) begin
      _T_1689 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1693 <= 22'h0;
    end else if (_T_1691) begin
      _T_1693 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1697 <= 22'h0;
    end else if (_T_1695) begin
      _T_1697 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1701 <= 22'h0;
    end else if (_T_1699) begin
      _T_1701 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1705 <= 22'h0;
    end else if (_T_1703) begin
      _T_1705 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1709 <= 22'h0;
    end else if (_T_1707) begin
      _T_1709 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1713 <= 22'h0;
    end else if (_T_1711) begin
      _T_1713 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1717 <= 22'h0;
    end else if (_T_1715) begin
      _T_1717 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1721 <= 22'h0;
    end else if (_T_1719) begin
      _T_1721 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1725 <= 22'h0;
    end else if (_T_1723) begin
      _T_1725 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1729 <= 22'h0;
    end else if (_T_1727) begin
      _T_1729 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1733 <= 22'h0;
    end else if (_T_1731) begin
      _T_1733 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1737 <= 22'h0;
    end else if (_T_1735) begin
      _T_1737 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1741 <= 22'h0;
    end else if (_T_1739) begin
      _T_1741 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1745 <= 22'h0;
    end else if (_T_1743) begin
      _T_1745 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1749 <= 22'h0;
    end else if (_T_1747) begin
      _T_1749 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1753 <= 22'h0;
    end else if (_T_1751) begin
      _T_1753 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1757 <= 22'h0;
    end else if (_T_1755) begin
      _T_1757 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1761 <= 22'h0;
    end else if (_T_1759) begin
      _T_1761 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1765 <= 22'h0;
    end else if (_T_1763) begin
      _T_1765 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1769 <= 22'h0;
    end else if (_T_1767) begin
      _T_1769 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1773 <= 22'h0;
    end else if (_T_1771) begin
      _T_1773 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1777 <= 22'h0;
    end else if (_T_1775) begin
      _T_1777 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1781 <= 22'h0;
    end else if (_T_1779) begin
      _T_1781 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1785 <= 22'h0;
    end else if (_T_1783) begin
      _T_1785 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1789 <= 22'h0;
    end else if (_T_1787) begin
      _T_1789 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1793 <= 22'h0;
    end else if (_T_1791) begin
      _T_1793 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1797 <= 22'h0;
    end else if (_T_1795) begin
      _T_1797 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1801 <= 22'h0;
    end else if (_T_1799) begin
      _T_1801 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1805 <= 22'h0;
    end else if (_T_1803) begin
      _T_1805 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1809 <= 22'h0;
    end else if (_T_1807) begin
      _T_1809 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1813 <= 22'h0;
    end else if (_T_1811) begin
      _T_1813 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1817 <= 22'h0;
    end else if (_T_1815) begin
      _T_1817 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1821 <= 22'h0;
    end else if (_T_1819) begin
      _T_1821 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1825 <= 22'h0;
    end else if (_T_1823) begin
      _T_1825 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1829 <= 22'h0;
    end else if (_T_1827) begin
      _T_1829 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1833 <= 22'h0;
    end else if (_T_1831) begin
      _T_1833 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1837 <= 22'h0;
    end else if (_T_1835) begin
      _T_1837 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1841 <= 22'h0;
    end else if (_T_1839) begin
      _T_1841 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1845 <= 22'h0;
    end else if (_T_1843) begin
      _T_1845 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1849 <= 22'h0;
    end else if (_T_1847) begin
      _T_1849 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1853 <= 22'h0;
    end else if (_T_1851) begin
      _T_1853 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1857 <= 22'h0;
    end else if (_T_1855) begin
      _T_1857 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1861 <= 22'h0;
    end else if (_T_1859) begin
      _T_1861 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1865 <= 22'h0;
    end else if (_T_1863) begin
      _T_1865 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1869 <= 22'h0;
    end else if (_T_1867) begin
      _T_1869 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1873 <= 22'h0;
    end else if (_T_1871) begin
      _T_1873 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1877 <= 22'h0;
    end else if (_T_1875) begin
      _T_1877 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1881 <= 22'h0;
    end else if (_T_1879) begin
      _T_1881 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1885 <= 22'h0;
    end else if (_T_1883) begin
      _T_1885 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1889 <= 22'h0;
    end else if (_T_1887) begin
      _T_1889 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1893 <= 22'h0;
    end else if (_T_1891) begin
      _T_1893 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1897 <= 22'h0;
    end else if (_T_1895) begin
      _T_1897 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1901 <= 22'h0;
    end else if (_T_1899) begin
      _T_1901 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1905 <= 22'h0;
    end else if (_T_1903) begin
      _T_1905 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1909 <= 22'h0;
    end else if (_T_1907) begin
      _T_1909 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1913 <= 22'h0;
    end else if (_T_1911) begin
      _T_1913 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1917 <= 22'h0;
    end else if (_T_1915) begin
      _T_1917 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1921 <= 22'h0;
    end else if (_T_1919) begin
      _T_1921 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1925 <= 22'h0;
    end else if (_T_1923) begin
      _T_1925 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1929 <= 22'h0;
    end else if (_T_1927) begin
      _T_1929 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1933 <= 22'h0;
    end else if (_T_1931) begin
      _T_1933 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1937 <= 22'h0;
    end else if (_T_1935) begin
      _T_1937 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1941 <= 22'h0;
    end else if (_T_1939) begin
      _T_1941 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1945 <= 22'h0;
    end else if (_T_1943) begin
      _T_1945 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1949 <= 22'h0;
    end else if (_T_1947) begin
      _T_1949 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1953 <= 22'h0;
    end else if (_T_1951) begin
      _T_1953 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1957 <= 22'h0;
    end else if (_T_1955) begin
      _T_1957 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1961 <= 22'h0;
    end else if (_T_1959) begin
      _T_1961 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1965 <= 22'h0;
    end else if (_T_1963) begin
      _T_1965 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1969 <= 22'h0;
    end else if (_T_1967) begin
      _T_1969 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1973 <= 22'h0;
    end else if (_T_1971) begin
      _T_1973 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1977 <= 22'h0;
    end else if (_T_1975) begin
      _T_1977 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1981 <= 22'h0;
    end else if (_T_1979) begin
      _T_1981 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1985 <= 22'h0;
    end else if (_T_1983) begin
      _T_1985 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1989 <= 22'h0;
    end else if (_T_1987) begin
      _T_1989 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1993 <= 22'h0;
    end else if (_T_1991) begin
      _T_1993 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1997 <= 22'h0;
    end else if (_T_1995) begin
      _T_1997 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2001 <= 22'h0;
    end else if (_T_1999) begin
      _T_2001 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2005 <= 22'h0;
    end else if (_T_2003) begin
      _T_2005 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2009 <= 22'h0;
    end else if (_T_2007) begin
      _T_2009 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2013 <= 22'h0;
    end else if (_T_2011) begin
      _T_2013 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2017 <= 22'h0;
    end else if (_T_2015) begin
      _T_2017 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2021 <= 22'h0;
    end else if (_T_2019) begin
      _T_2021 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2025 <= 22'h0;
    end else if (_T_2023) begin
      _T_2025 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2029 <= 22'h0;
    end else if (_T_2027) begin
      _T_2029 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2033 <= 22'h0;
    end else if (_T_2031) begin
      _T_2033 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2037 <= 22'h0;
    end else if (_T_2035) begin
      _T_2037 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2041 <= 22'h0;
    end else if (_T_2039) begin
      _T_2041 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2045 <= 22'h0;
    end else if (_T_2043) begin
      _T_2045 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2049 <= 22'h0;
    end else if (_T_2047) begin
      _T_2049 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2053 <= 22'h0;
    end else if (_T_2051) begin
      _T_2053 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2057 <= 22'h0;
    end else if (_T_2055) begin
      _T_2057 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2061 <= 22'h0;
    end else if (_T_2059) begin
      _T_2061 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2065 <= 22'h0;
    end else if (_T_2063) begin
      _T_2065 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2069 <= 22'h0;
    end else if (_T_2067) begin
      _T_2069 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2073 <= 22'h0;
    end else if (_T_2071) begin
      _T_2073 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2077 <= 22'h0;
    end else if (_T_2075) begin
      _T_2077 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2081 <= 22'h0;
    end else if (_T_2079) begin
      _T_2081 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2085 <= 22'h0;
    end else if (_T_2083) begin
      _T_2085 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2089 <= 22'h0;
    end else if (_T_2087) begin
      _T_2089 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2093 <= 22'h0;
    end else if (_T_2091) begin
      _T_2093 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2097 <= 22'h0;
    end else if (_T_2095) begin
      _T_2097 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2101 <= 22'h0;
    end else if (_T_2099) begin
      _T_2101 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2105 <= 22'h0;
    end else if (_T_2103) begin
      _T_2105 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2109 <= 22'h0;
    end else if (_T_2107) begin
      _T_2109 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2113 <= 22'h0;
    end else if (_T_2111) begin
      _T_2113 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2117 <= 22'h0;
    end else if (_T_2115) begin
      _T_2117 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2121 <= 22'h0;
    end else if (_T_2119) begin
      _T_2121 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2125 <= 22'h0;
    end else if (_T_2123) begin
      _T_2125 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2129 <= 22'h0;
    end else if (_T_2127) begin
      _T_2129 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2133 <= 22'h0;
    end else if (_T_2131) begin
      _T_2133 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2137 <= 22'h0;
    end else if (_T_2135) begin
      _T_2137 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2141 <= 22'h0;
    end else if (_T_2139) begin
      _T_2141 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2145 <= 22'h0;
    end else if (_T_2143) begin
      _T_2145 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2149 <= 22'h0;
    end else if (_T_2147) begin
      _T_2149 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2153 <= 22'h0;
    end else if (_T_2151) begin
      _T_2153 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2157 <= 22'h0;
    end else if (_T_2155) begin
      _T_2157 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2161 <= 22'h0;
    end else if (_T_2159) begin
      _T_2161 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2165 <= 22'h0;
    end else if (_T_2163) begin
      _T_2165 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2169 <= 22'h0;
    end else if (_T_2167) begin
      _T_2169 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2173 <= 22'h0;
    end else if (_T_2171) begin
      _T_2173 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2177 <= 22'h0;
    end else if (_T_2175) begin
      _T_2177 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2181 <= 22'h0;
    end else if (_T_2179) begin
      _T_2181 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2185 <= 22'h0;
    end else if (_T_2183) begin
      _T_2185 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2189 <= 22'h0;
    end else if (_T_2187) begin
      _T_2189 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2193 <= 22'h0;
    end else if (_T_2191) begin
      _T_2193 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2197 <= 22'h0;
    end else if (_T_2195) begin
      _T_2197 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2201 <= 22'h0;
    end else if (_T_2199) begin
      _T_2201 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2205 <= 22'h0;
    end else if (_T_2203) begin
      _T_2205 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2209 <= 22'h0;
    end else if (_T_2207) begin
      _T_2209 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2213 <= 22'h0;
    end else if (_T_2211) begin
      _T_2213 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2217 <= 22'h0;
    end else if (_T_2215) begin
      _T_2217 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2221 <= 22'h0;
    end else if (_T_2219) begin
      _T_2221 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2225 <= 22'h0;
    end else if (_T_2223) begin
      _T_2225 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2229 <= 22'h0;
    end else if (_T_2227) begin
      _T_2229 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2233 <= 22'h0;
    end else if (_T_2231) begin
      _T_2233 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2237 <= 22'h0;
    end else if (_T_2235) begin
      _T_2237 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2241 <= 22'h0;
    end else if (_T_2239) begin
      _T_2241 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2245 <= 22'h0;
    end else if (_T_2243) begin
      _T_2245 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2249 <= 22'h0;
    end else if (_T_2247) begin
      _T_2249 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2253 <= 22'h0;
    end else if (_T_2251) begin
      _T_2253 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2257 <= 22'h0;
    end else if (_T_2255) begin
      _T_2257 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2261 <= 22'h0;
    end else if (_T_2259) begin
      _T_2261 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2265 <= 22'h0;
    end else if (_T_2263) begin
      _T_2265 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2269 <= 22'h0;
    end else if (_T_2267) begin
      _T_2269 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2273 <= 22'h0;
    end else if (_T_2271) begin
      _T_2273 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2277 <= 22'h0;
    end else if (_T_2275) begin
      _T_2277 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2281 <= 22'h0;
    end else if (_T_2279) begin
      _T_2281 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2285 <= 22'h0;
    end else if (_T_2283) begin
      _T_2285 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2289 <= 22'h0;
    end else if (_T_2287) begin
      _T_2289 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2293 <= 22'h0;
    end else if (_T_2291) begin
      _T_2293 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2297 <= 22'h0;
    end else if (_T_2295) begin
      _T_2297 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2301 <= 22'h0;
    end else if (_T_2299) begin
      _T_2301 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2305 <= 22'h0;
    end else if (_T_2303) begin
      _T_2305 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2309 <= 22'h0;
    end else if (_T_2307) begin
      _T_2309 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2313 <= 22'h0;
    end else if (_T_2311) begin
      _T_2313 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2317 <= 22'h0;
    end else if (_T_2315) begin
      _T_2317 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2321 <= 22'h0;
    end else if (_T_2319) begin
      _T_2321 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2325 <= 22'h0;
    end else if (_T_2323) begin
      _T_2325 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2329 <= 22'h0;
    end else if (_T_2327) begin
      _T_2329 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2333 <= 22'h0;
    end else if (_T_2331) begin
      _T_2333 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2337 <= 22'h0;
    end else if (_T_2335) begin
      _T_2337 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2341 <= 22'h0;
    end else if (_T_2339) begin
      _T_2341 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2345 <= 22'h0;
    end else if (_T_2343) begin
      _T_2345 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2349 <= 22'h0;
    end else if (_T_2347) begin
      _T_2349 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2353 <= 22'h0;
    end else if (_T_2351) begin
      _T_2353 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2357 <= 22'h0;
    end else if (_T_2355) begin
      _T_2357 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2361 <= 22'h0;
    end else if (_T_2359) begin
      _T_2361 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2365 <= 22'h0;
    end else if (_T_2363) begin
      _T_2365 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2369 <= 22'h0;
    end else if (_T_2367) begin
      _T_2369 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2373 <= 22'h0;
    end else if (_T_2371) begin
      _T_2373 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2377 <= 22'h0;
    end else if (_T_2375) begin
      _T_2377 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2381 <= 22'h0;
    end else if (_T_2379) begin
      _T_2381 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2385 <= 22'h0;
    end else if (_T_2383) begin
      _T_2385 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2389 <= 22'h0;
    end else if (_T_2387) begin
      _T_2389 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2393 <= 22'h0;
    end else if (_T_2391) begin
      _T_2393 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2397 <= 22'h0;
    end else if (_T_2395) begin
      _T_2397 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2401 <= 22'h0;
    end else if (_T_2399) begin
      _T_2401 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2405 <= 22'h0;
    end else if (_T_2403) begin
      _T_2405 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2409 <= 22'h0;
    end else if (_T_2407) begin
      _T_2409 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2413 <= 22'h0;
    end else if (_T_2411) begin
      _T_2413 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2417 <= 22'h0;
    end else if (_T_2415) begin
      _T_2417 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2421 <= 22'h0;
    end else if (_T_2419) begin
      _T_2421 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2425 <= 22'h0;
    end else if (_T_2423) begin
      _T_2425 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2429 <= 22'h0;
    end else if (_T_2427) begin
      _T_2429 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2433 <= 22'h0;
    end else if (_T_2431) begin
      _T_2433 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2437 <= 22'h0;
    end else if (_T_2435) begin
      _T_2437 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2441 <= 22'h0;
    end else if (_T_2439) begin
      _T_2441 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2445 <= 22'h0;
    end else if (_T_2443) begin
      _T_2445 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2449 <= 22'h0;
    end else if (_T_2447) begin
      _T_2449 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2453 <= 22'h0;
    end else if (_T_2451) begin
      _T_2453 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2457 <= 22'h0;
    end else if (_T_2455) begin
      _T_2457 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2461 <= 22'h0;
    end else if (_T_2459) begin
      _T_2461 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2465 <= 22'h0;
    end else if (_T_2463) begin
      _T_2465 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2469 <= 22'h0;
    end else if (_T_2467) begin
      _T_2469 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2473 <= 22'h0;
    end else if (_T_2471) begin
      _T_2473 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2477 <= 22'h0;
    end else if (_T_2475) begin
      _T_2477 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2481 <= 22'h0;
    end else if (_T_2479) begin
      _T_2481 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2485 <= 22'h0;
    end else if (_T_2483) begin
      _T_2485 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2489 <= 22'h0;
    end else if (_T_2487) begin
      _T_2489 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2493 <= 22'h0;
    end else if (_T_2491) begin
      _T_2493 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2497 <= 22'h0;
    end else if (_T_2495) begin
      _T_2497 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2501 <= 22'h0;
    end else if (_T_2499) begin
      _T_2501 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2505 <= 22'h0;
    end else if (_T_2503) begin
      _T_2505 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2509 <= 22'h0;
    end else if (_T_2507) begin
      _T_2509 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2513 <= 22'h0;
    end else if (_T_2511) begin
      _T_2513 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2517 <= 22'h0;
    end else if (_T_2515) begin
      _T_2517 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2521 <= 22'h0;
    end else if (_T_2519) begin
      _T_2521 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2525 <= 22'h0;
    end else if (_T_2523) begin
      _T_2525 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2529 <= 22'h0;
    end else if (_T_2527) begin
      _T_2529 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2533 <= 22'h0;
    end else if (_T_2531) begin
      _T_2533 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2537 <= 22'h0;
    end else if (_T_2535) begin
      _T_2537 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2541 <= 22'h0;
    end else if (_T_2539) begin
      _T_2541 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2545 <= 22'h0;
    end else if (_T_2543) begin
      _T_2545 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2549 <= 22'h0;
    end else if (_T_2547) begin
      _T_2549 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2553 <= 22'h0;
    end else if (_T_2551) begin
      _T_2553 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2557 <= 22'h0;
    end else if (_T_2555) begin
      _T_2557 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2561 <= 22'h0;
    end else if (_T_2559) begin
      _T_2561 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2565 <= 22'h0;
    end else if (_T_2563) begin
      _T_2565 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2569 <= 22'h0;
    end else if (_T_2567) begin
      _T_2569 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2573 <= 22'h0;
    end else if (_T_2571) begin
      _T_2573 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2577 <= 22'h0;
    end else if (_T_2575) begin
      _T_2577 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2581 <= 22'h0;
    end else if (_T_2579) begin
      _T_2581 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2585 <= 22'h0;
    end else if (_T_2583) begin
      _T_2585 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2589 <= 22'h0;
    end else if (_T_2587) begin
      _T_2589 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2593 <= 22'h0;
    end else if (_T_2591) begin
      _T_2593 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2597 <= 22'h0;
    end else if (_T_2595) begin
      _T_2597 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2601 <= 22'h0;
    end else if (_T_2599) begin
      _T_2601 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2605 <= 22'h0;
    end else if (_T_2603) begin
      _T_2605 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2609 <= 22'h0;
    end else if (_T_2607) begin
      _T_2609 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2613 <= 22'h0;
    end else if (_T_2611) begin
      _T_2613 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2617 <= 22'h0;
    end else if (_T_2615) begin
      _T_2617 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2621 <= 22'h0;
    end else if (_T_2619) begin
      _T_2621 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2625 <= 22'h0;
    end else if (_T_2623) begin
      _T_2625 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2629 <= 22'h0;
    end else if (_T_2627) begin
      _T_2629 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2633 <= 22'h0;
    end else if (_T_2631) begin
      _T_2633 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2637 <= 22'h0;
    end else if (_T_2635) begin
      _T_2637 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2641 <= 22'h0;
    end else if (_T_2639) begin
      _T_2641 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2645 <= 22'h0;
    end else if (_T_2643) begin
      _T_2645 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2649 <= 22'h0;
    end else if (_T_2647) begin
      _T_2649 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2653 <= 22'h0;
    end else if (_T_2651) begin
      _T_2653 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2657 <= 22'h0;
    end else if (_T_2655) begin
      _T_2657 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2661 <= 22'h0;
    end else if (_T_2659) begin
      _T_2661 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2665 <= 22'h0;
    end else if (_T_2663) begin
      _T_2665 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2669 <= 22'h0;
    end else if (_T_2667) begin
      _T_2669 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2673 <= 22'h0;
    end else if (_T_2671) begin
      _T_2673 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2677 <= 22'h0;
    end else if (_T_2675) begin
      _T_2677 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2681 <= 22'h0;
    end else if (_T_2679) begin
      _T_2681 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2685 <= 22'h0;
    end else if (_T_2683) begin
      _T_2685 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_2689 <= 22'h0;
    end else if (_T_2687) begin
      _T_2689 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      fghr <= 8'h0;
    end else if (_T_375) begin
      fghr <= fghr_ns;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_0 <= 2'h0;
    end else if (bht_bank_sel_1_0_0) begin
      if (_T_9449) begin
        bht_bank_rd_data_out_1_0 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_0 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_1 <= 2'h0;
    end else if (bht_bank_sel_1_0_1) begin
      if (_T_9458) begin
        bht_bank_rd_data_out_1_1 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_1 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_2 <= 2'h0;
    end else if (bht_bank_sel_1_0_2) begin
      if (_T_9467) begin
        bht_bank_rd_data_out_1_2 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_2 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_3 <= 2'h0;
    end else if (bht_bank_sel_1_0_3) begin
      if (_T_9476) begin
        bht_bank_rd_data_out_1_3 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_3 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_4 <= 2'h0;
    end else if (bht_bank_sel_1_0_4) begin
      if (_T_9485) begin
        bht_bank_rd_data_out_1_4 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_4 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_5 <= 2'h0;
    end else if (bht_bank_sel_1_0_5) begin
      if (_T_9494) begin
        bht_bank_rd_data_out_1_5 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_5 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_6 <= 2'h0;
    end else if (bht_bank_sel_1_0_6) begin
      if (_T_9503) begin
        bht_bank_rd_data_out_1_6 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_6 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_7 <= 2'h0;
    end else if (bht_bank_sel_1_0_7) begin
      if (_T_9512) begin
        bht_bank_rd_data_out_1_7 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_7 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_8 <= 2'h0;
    end else if (bht_bank_sel_1_0_8) begin
      if (_T_9521) begin
        bht_bank_rd_data_out_1_8 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_8 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_9 <= 2'h0;
    end else if (bht_bank_sel_1_0_9) begin
      if (_T_9530) begin
        bht_bank_rd_data_out_1_9 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_9 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_10 <= 2'h0;
    end else if (bht_bank_sel_1_0_10) begin
      if (_T_9539) begin
        bht_bank_rd_data_out_1_10 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_10 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_11 <= 2'h0;
    end else if (bht_bank_sel_1_0_11) begin
      if (_T_9548) begin
        bht_bank_rd_data_out_1_11 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_11 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_12 <= 2'h0;
    end else if (bht_bank_sel_1_0_12) begin
      if (_T_9557) begin
        bht_bank_rd_data_out_1_12 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_12 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_13 <= 2'h0;
    end else if (bht_bank_sel_1_0_13) begin
      if (_T_9566) begin
        bht_bank_rd_data_out_1_13 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_13 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_14 <= 2'h0;
    end else if (bht_bank_sel_1_0_14) begin
      if (_T_9575) begin
        bht_bank_rd_data_out_1_14 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_14 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_15 <= 2'h0;
    end else if (bht_bank_sel_1_0_15) begin
      if (_T_9584) begin
        bht_bank_rd_data_out_1_15 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_15 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_16 <= 2'h0;
    end else if (bht_bank_sel_1_1_0) begin
      if (_T_9593) begin
        bht_bank_rd_data_out_1_16 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_16 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_17 <= 2'h0;
    end else if (bht_bank_sel_1_1_1) begin
      if (_T_9602) begin
        bht_bank_rd_data_out_1_17 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_17 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_18 <= 2'h0;
    end else if (bht_bank_sel_1_1_2) begin
      if (_T_9611) begin
        bht_bank_rd_data_out_1_18 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_18 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_19 <= 2'h0;
    end else if (bht_bank_sel_1_1_3) begin
      if (_T_9620) begin
        bht_bank_rd_data_out_1_19 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_19 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_20 <= 2'h0;
    end else if (bht_bank_sel_1_1_4) begin
      if (_T_9629) begin
        bht_bank_rd_data_out_1_20 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_20 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_21 <= 2'h0;
    end else if (bht_bank_sel_1_1_5) begin
      if (_T_9638) begin
        bht_bank_rd_data_out_1_21 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_21 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_22 <= 2'h0;
    end else if (bht_bank_sel_1_1_6) begin
      if (_T_9647) begin
        bht_bank_rd_data_out_1_22 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_22 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_23 <= 2'h0;
    end else if (bht_bank_sel_1_1_7) begin
      if (_T_9656) begin
        bht_bank_rd_data_out_1_23 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_23 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_24 <= 2'h0;
    end else if (bht_bank_sel_1_1_8) begin
      if (_T_9665) begin
        bht_bank_rd_data_out_1_24 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_24 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_25 <= 2'h0;
    end else if (bht_bank_sel_1_1_9) begin
      if (_T_9674) begin
        bht_bank_rd_data_out_1_25 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_25 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_26 <= 2'h0;
    end else if (bht_bank_sel_1_1_10) begin
      if (_T_9683) begin
        bht_bank_rd_data_out_1_26 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_26 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_27 <= 2'h0;
    end else if (bht_bank_sel_1_1_11) begin
      if (_T_9692) begin
        bht_bank_rd_data_out_1_27 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_27 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_28 <= 2'h0;
    end else if (bht_bank_sel_1_1_12) begin
      if (_T_9701) begin
        bht_bank_rd_data_out_1_28 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_28 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_29 <= 2'h0;
    end else if (bht_bank_sel_1_1_13) begin
      if (_T_9710) begin
        bht_bank_rd_data_out_1_29 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_29 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_30 <= 2'h0;
    end else if (bht_bank_sel_1_1_14) begin
      if (_T_9719) begin
        bht_bank_rd_data_out_1_30 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_30 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_31 <= 2'h0;
    end else if (bht_bank_sel_1_1_15) begin
      if (_T_9728) begin
        bht_bank_rd_data_out_1_31 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_31 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_32 <= 2'h0;
    end else if (bht_bank_sel_1_2_0) begin
      if (_T_9737) begin
        bht_bank_rd_data_out_1_32 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_32 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_33 <= 2'h0;
    end else if (bht_bank_sel_1_2_1) begin
      if (_T_9746) begin
        bht_bank_rd_data_out_1_33 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_33 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_34 <= 2'h0;
    end else if (bht_bank_sel_1_2_2) begin
      if (_T_9755) begin
        bht_bank_rd_data_out_1_34 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_34 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_35 <= 2'h0;
    end else if (bht_bank_sel_1_2_3) begin
      if (_T_9764) begin
        bht_bank_rd_data_out_1_35 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_35 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_36 <= 2'h0;
    end else if (bht_bank_sel_1_2_4) begin
      if (_T_9773) begin
        bht_bank_rd_data_out_1_36 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_36 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_37 <= 2'h0;
    end else if (bht_bank_sel_1_2_5) begin
      if (_T_9782) begin
        bht_bank_rd_data_out_1_37 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_37 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_38 <= 2'h0;
    end else if (bht_bank_sel_1_2_6) begin
      if (_T_9791) begin
        bht_bank_rd_data_out_1_38 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_38 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_39 <= 2'h0;
    end else if (bht_bank_sel_1_2_7) begin
      if (_T_9800) begin
        bht_bank_rd_data_out_1_39 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_39 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_40 <= 2'h0;
    end else if (bht_bank_sel_1_2_8) begin
      if (_T_9809) begin
        bht_bank_rd_data_out_1_40 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_40 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_41 <= 2'h0;
    end else if (bht_bank_sel_1_2_9) begin
      if (_T_9818) begin
        bht_bank_rd_data_out_1_41 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_41 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_42 <= 2'h0;
    end else if (bht_bank_sel_1_2_10) begin
      if (_T_9827) begin
        bht_bank_rd_data_out_1_42 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_42 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_43 <= 2'h0;
    end else if (bht_bank_sel_1_2_11) begin
      if (_T_9836) begin
        bht_bank_rd_data_out_1_43 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_43 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_44 <= 2'h0;
    end else if (bht_bank_sel_1_2_12) begin
      if (_T_9845) begin
        bht_bank_rd_data_out_1_44 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_44 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_45 <= 2'h0;
    end else if (bht_bank_sel_1_2_13) begin
      if (_T_9854) begin
        bht_bank_rd_data_out_1_45 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_45 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_46 <= 2'h0;
    end else if (bht_bank_sel_1_2_14) begin
      if (_T_9863) begin
        bht_bank_rd_data_out_1_46 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_46 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_47 <= 2'h0;
    end else if (bht_bank_sel_1_2_15) begin
      if (_T_9872) begin
        bht_bank_rd_data_out_1_47 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_47 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_48 <= 2'h0;
    end else if (bht_bank_sel_1_3_0) begin
      if (_T_9881) begin
        bht_bank_rd_data_out_1_48 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_48 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_49 <= 2'h0;
    end else if (bht_bank_sel_1_3_1) begin
      if (_T_9890) begin
        bht_bank_rd_data_out_1_49 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_49 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_50 <= 2'h0;
    end else if (bht_bank_sel_1_3_2) begin
      if (_T_9899) begin
        bht_bank_rd_data_out_1_50 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_50 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_51 <= 2'h0;
    end else if (bht_bank_sel_1_3_3) begin
      if (_T_9908) begin
        bht_bank_rd_data_out_1_51 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_51 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_52 <= 2'h0;
    end else if (bht_bank_sel_1_3_4) begin
      if (_T_9917) begin
        bht_bank_rd_data_out_1_52 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_52 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_53 <= 2'h0;
    end else if (bht_bank_sel_1_3_5) begin
      if (_T_9926) begin
        bht_bank_rd_data_out_1_53 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_53 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_54 <= 2'h0;
    end else if (bht_bank_sel_1_3_6) begin
      if (_T_9935) begin
        bht_bank_rd_data_out_1_54 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_54 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_55 <= 2'h0;
    end else if (bht_bank_sel_1_3_7) begin
      if (_T_9944) begin
        bht_bank_rd_data_out_1_55 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_55 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_56 <= 2'h0;
    end else if (bht_bank_sel_1_3_8) begin
      if (_T_9953) begin
        bht_bank_rd_data_out_1_56 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_56 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_57 <= 2'h0;
    end else if (bht_bank_sel_1_3_9) begin
      if (_T_9962) begin
        bht_bank_rd_data_out_1_57 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_57 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_58 <= 2'h0;
    end else if (bht_bank_sel_1_3_10) begin
      if (_T_9971) begin
        bht_bank_rd_data_out_1_58 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_58 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_59 <= 2'h0;
    end else if (bht_bank_sel_1_3_11) begin
      if (_T_9980) begin
        bht_bank_rd_data_out_1_59 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_59 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_60 <= 2'h0;
    end else if (bht_bank_sel_1_3_12) begin
      if (_T_9989) begin
        bht_bank_rd_data_out_1_60 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_60 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_61 <= 2'h0;
    end else if (bht_bank_sel_1_3_13) begin
      if (_T_9998) begin
        bht_bank_rd_data_out_1_61 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_61 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_62 <= 2'h0;
    end else if (bht_bank_sel_1_3_14) begin
      if (_T_10007) begin
        bht_bank_rd_data_out_1_62 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_62 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_63 <= 2'h0;
    end else if (bht_bank_sel_1_3_15) begin
      if (_T_10016) begin
        bht_bank_rd_data_out_1_63 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_63 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_64 <= 2'h0;
    end else if (bht_bank_sel_1_4_0) begin
      if (_T_10025) begin
        bht_bank_rd_data_out_1_64 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_64 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_65 <= 2'h0;
    end else if (bht_bank_sel_1_4_1) begin
      if (_T_10034) begin
        bht_bank_rd_data_out_1_65 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_65 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_66 <= 2'h0;
    end else if (bht_bank_sel_1_4_2) begin
      if (_T_10043) begin
        bht_bank_rd_data_out_1_66 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_66 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_67 <= 2'h0;
    end else if (bht_bank_sel_1_4_3) begin
      if (_T_10052) begin
        bht_bank_rd_data_out_1_67 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_67 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_68 <= 2'h0;
    end else if (bht_bank_sel_1_4_4) begin
      if (_T_10061) begin
        bht_bank_rd_data_out_1_68 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_68 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_69 <= 2'h0;
    end else if (bht_bank_sel_1_4_5) begin
      if (_T_10070) begin
        bht_bank_rd_data_out_1_69 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_69 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_70 <= 2'h0;
    end else if (bht_bank_sel_1_4_6) begin
      if (_T_10079) begin
        bht_bank_rd_data_out_1_70 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_70 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_71 <= 2'h0;
    end else if (bht_bank_sel_1_4_7) begin
      if (_T_10088) begin
        bht_bank_rd_data_out_1_71 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_71 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_72 <= 2'h0;
    end else if (bht_bank_sel_1_4_8) begin
      if (_T_10097) begin
        bht_bank_rd_data_out_1_72 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_72 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_73 <= 2'h0;
    end else if (bht_bank_sel_1_4_9) begin
      if (_T_10106) begin
        bht_bank_rd_data_out_1_73 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_73 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_74 <= 2'h0;
    end else if (bht_bank_sel_1_4_10) begin
      if (_T_10115) begin
        bht_bank_rd_data_out_1_74 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_74 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_75 <= 2'h0;
    end else if (bht_bank_sel_1_4_11) begin
      if (_T_10124) begin
        bht_bank_rd_data_out_1_75 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_75 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_76 <= 2'h0;
    end else if (bht_bank_sel_1_4_12) begin
      if (_T_10133) begin
        bht_bank_rd_data_out_1_76 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_76 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_77 <= 2'h0;
    end else if (bht_bank_sel_1_4_13) begin
      if (_T_10142) begin
        bht_bank_rd_data_out_1_77 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_77 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_78 <= 2'h0;
    end else if (bht_bank_sel_1_4_14) begin
      if (_T_10151) begin
        bht_bank_rd_data_out_1_78 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_78 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_79 <= 2'h0;
    end else if (bht_bank_sel_1_4_15) begin
      if (_T_10160) begin
        bht_bank_rd_data_out_1_79 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_79 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_80 <= 2'h0;
    end else if (bht_bank_sel_1_5_0) begin
      if (_T_10169) begin
        bht_bank_rd_data_out_1_80 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_80 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_81 <= 2'h0;
    end else if (bht_bank_sel_1_5_1) begin
      if (_T_10178) begin
        bht_bank_rd_data_out_1_81 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_81 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_82 <= 2'h0;
    end else if (bht_bank_sel_1_5_2) begin
      if (_T_10187) begin
        bht_bank_rd_data_out_1_82 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_82 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_83 <= 2'h0;
    end else if (bht_bank_sel_1_5_3) begin
      if (_T_10196) begin
        bht_bank_rd_data_out_1_83 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_83 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_84 <= 2'h0;
    end else if (bht_bank_sel_1_5_4) begin
      if (_T_10205) begin
        bht_bank_rd_data_out_1_84 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_84 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_85 <= 2'h0;
    end else if (bht_bank_sel_1_5_5) begin
      if (_T_10214) begin
        bht_bank_rd_data_out_1_85 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_85 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_86 <= 2'h0;
    end else if (bht_bank_sel_1_5_6) begin
      if (_T_10223) begin
        bht_bank_rd_data_out_1_86 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_86 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_87 <= 2'h0;
    end else if (bht_bank_sel_1_5_7) begin
      if (_T_10232) begin
        bht_bank_rd_data_out_1_87 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_87 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_88 <= 2'h0;
    end else if (bht_bank_sel_1_5_8) begin
      if (_T_10241) begin
        bht_bank_rd_data_out_1_88 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_88 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_89 <= 2'h0;
    end else if (bht_bank_sel_1_5_9) begin
      if (_T_10250) begin
        bht_bank_rd_data_out_1_89 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_89 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_90 <= 2'h0;
    end else if (bht_bank_sel_1_5_10) begin
      if (_T_10259) begin
        bht_bank_rd_data_out_1_90 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_90 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_91 <= 2'h0;
    end else if (bht_bank_sel_1_5_11) begin
      if (_T_10268) begin
        bht_bank_rd_data_out_1_91 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_91 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_92 <= 2'h0;
    end else if (bht_bank_sel_1_5_12) begin
      if (_T_10277) begin
        bht_bank_rd_data_out_1_92 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_92 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_93 <= 2'h0;
    end else if (bht_bank_sel_1_5_13) begin
      if (_T_10286) begin
        bht_bank_rd_data_out_1_93 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_93 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_94 <= 2'h0;
    end else if (bht_bank_sel_1_5_14) begin
      if (_T_10295) begin
        bht_bank_rd_data_out_1_94 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_94 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_95 <= 2'h0;
    end else if (bht_bank_sel_1_5_15) begin
      if (_T_10304) begin
        bht_bank_rd_data_out_1_95 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_95 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_96 <= 2'h0;
    end else if (bht_bank_sel_1_6_0) begin
      if (_T_10313) begin
        bht_bank_rd_data_out_1_96 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_96 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_97 <= 2'h0;
    end else if (bht_bank_sel_1_6_1) begin
      if (_T_10322) begin
        bht_bank_rd_data_out_1_97 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_97 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_98 <= 2'h0;
    end else if (bht_bank_sel_1_6_2) begin
      if (_T_10331) begin
        bht_bank_rd_data_out_1_98 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_98 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_99 <= 2'h0;
    end else if (bht_bank_sel_1_6_3) begin
      if (_T_10340) begin
        bht_bank_rd_data_out_1_99 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_99 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_100 <= 2'h0;
    end else if (bht_bank_sel_1_6_4) begin
      if (_T_10349) begin
        bht_bank_rd_data_out_1_100 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_100 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_101 <= 2'h0;
    end else if (bht_bank_sel_1_6_5) begin
      if (_T_10358) begin
        bht_bank_rd_data_out_1_101 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_101 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_102 <= 2'h0;
    end else if (bht_bank_sel_1_6_6) begin
      if (_T_10367) begin
        bht_bank_rd_data_out_1_102 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_102 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_103 <= 2'h0;
    end else if (bht_bank_sel_1_6_7) begin
      if (_T_10376) begin
        bht_bank_rd_data_out_1_103 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_103 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_104 <= 2'h0;
    end else if (bht_bank_sel_1_6_8) begin
      if (_T_10385) begin
        bht_bank_rd_data_out_1_104 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_104 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_105 <= 2'h0;
    end else if (bht_bank_sel_1_6_9) begin
      if (_T_10394) begin
        bht_bank_rd_data_out_1_105 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_105 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_106 <= 2'h0;
    end else if (bht_bank_sel_1_6_10) begin
      if (_T_10403) begin
        bht_bank_rd_data_out_1_106 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_106 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_107 <= 2'h0;
    end else if (bht_bank_sel_1_6_11) begin
      if (_T_10412) begin
        bht_bank_rd_data_out_1_107 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_107 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_108 <= 2'h0;
    end else if (bht_bank_sel_1_6_12) begin
      if (_T_10421) begin
        bht_bank_rd_data_out_1_108 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_108 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_109 <= 2'h0;
    end else if (bht_bank_sel_1_6_13) begin
      if (_T_10430) begin
        bht_bank_rd_data_out_1_109 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_109 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_110 <= 2'h0;
    end else if (bht_bank_sel_1_6_14) begin
      if (_T_10439) begin
        bht_bank_rd_data_out_1_110 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_110 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_111 <= 2'h0;
    end else if (bht_bank_sel_1_6_15) begin
      if (_T_10448) begin
        bht_bank_rd_data_out_1_111 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_111 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_112 <= 2'h0;
    end else if (bht_bank_sel_1_7_0) begin
      if (_T_10457) begin
        bht_bank_rd_data_out_1_112 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_112 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_113 <= 2'h0;
    end else if (bht_bank_sel_1_7_1) begin
      if (_T_10466) begin
        bht_bank_rd_data_out_1_113 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_113 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_114 <= 2'h0;
    end else if (bht_bank_sel_1_7_2) begin
      if (_T_10475) begin
        bht_bank_rd_data_out_1_114 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_114 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_115 <= 2'h0;
    end else if (bht_bank_sel_1_7_3) begin
      if (_T_10484) begin
        bht_bank_rd_data_out_1_115 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_115 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_116 <= 2'h0;
    end else if (bht_bank_sel_1_7_4) begin
      if (_T_10493) begin
        bht_bank_rd_data_out_1_116 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_116 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_117 <= 2'h0;
    end else if (bht_bank_sel_1_7_5) begin
      if (_T_10502) begin
        bht_bank_rd_data_out_1_117 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_117 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_118 <= 2'h0;
    end else if (bht_bank_sel_1_7_6) begin
      if (_T_10511) begin
        bht_bank_rd_data_out_1_118 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_118 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_119 <= 2'h0;
    end else if (bht_bank_sel_1_7_7) begin
      if (_T_10520) begin
        bht_bank_rd_data_out_1_119 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_119 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_120 <= 2'h0;
    end else if (bht_bank_sel_1_7_8) begin
      if (_T_10529) begin
        bht_bank_rd_data_out_1_120 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_120 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_121 <= 2'h0;
    end else if (bht_bank_sel_1_7_9) begin
      if (_T_10538) begin
        bht_bank_rd_data_out_1_121 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_121 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_122 <= 2'h0;
    end else if (bht_bank_sel_1_7_10) begin
      if (_T_10547) begin
        bht_bank_rd_data_out_1_122 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_122 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_123 <= 2'h0;
    end else if (bht_bank_sel_1_7_11) begin
      if (_T_10556) begin
        bht_bank_rd_data_out_1_123 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_123 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_124 <= 2'h0;
    end else if (bht_bank_sel_1_7_12) begin
      if (_T_10565) begin
        bht_bank_rd_data_out_1_124 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_124 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_125 <= 2'h0;
    end else if (bht_bank_sel_1_7_13) begin
      if (_T_10574) begin
        bht_bank_rd_data_out_1_125 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_125 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_126 <= 2'h0;
    end else if (bht_bank_sel_1_7_14) begin
      if (_T_10583) begin
        bht_bank_rd_data_out_1_126 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_126 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_127 <= 2'h0;
    end else if (bht_bank_sel_1_7_15) begin
      if (_T_10592) begin
        bht_bank_rd_data_out_1_127 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_127 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_128 <= 2'h0;
    end else if (bht_bank_sel_1_8_0) begin
      if (_T_10601) begin
        bht_bank_rd_data_out_1_128 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_128 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_129 <= 2'h0;
    end else if (bht_bank_sel_1_8_1) begin
      if (_T_10610) begin
        bht_bank_rd_data_out_1_129 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_129 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_130 <= 2'h0;
    end else if (bht_bank_sel_1_8_2) begin
      if (_T_10619) begin
        bht_bank_rd_data_out_1_130 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_130 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_131 <= 2'h0;
    end else if (bht_bank_sel_1_8_3) begin
      if (_T_10628) begin
        bht_bank_rd_data_out_1_131 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_131 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_132 <= 2'h0;
    end else if (bht_bank_sel_1_8_4) begin
      if (_T_10637) begin
        bht_bank_rd_data_out_1_132 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_132 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_133 <= 2'h0;
    end else if (bht_bank_sel_1_8_5) begin
      if (_T_10646) begin
        bht_bank_rd_data_out_1_133 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_133 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_134 <= 2'h0;
    end else if (bht_bank_sel_1_8_6) begin
      if (_T_10655) begin
        bht_bank_rd_data_out_1_134 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_134 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_135 <= 2'h0;
    end else if (bht_bank_sel_1_8_7) begin
      if (_T_10664) begin
        bht_bank_rd_data_out_1_135 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_135 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_136 <= 2'h0;
    end else if (bht_bank_sel_1_8_8) begin
      if (_T_10673) begin
        bht_bank_rd_data_out_1_136 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_136 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_137 <= 2'h0;
    end else if (bht_bank_sel_1_8_9) begin
      if (_T_10682) begin
        bht_bank_rd_data_out_1_137 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_137 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_138 <= 2'h0;
    end else if (bht_bank_sel_1_8_10) begin
      if (_T_10691) begin
        bht_bank_rd_data_out_1_138 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_138 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_139 <= 2'h0;
    end else if (bht_bank_sel_1_8_11) begin
      if (_T_10700) begin
        bht_bank_rd_data_out_1_139 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_139 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_140 <= 2'h0;
    end else if (bht_bank_sel_1_8_12) begin
      if (_T_10709) begin
        bht_bank_rd_data_out_1_140 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_140 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_141 <= 2'h0;
    end else if (bht_bank_sel_1_8_13) begin
      if (_T_10718) begin
        bht_bank_rd_data_out_1_141 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_141 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_142 <= 2'h0;
    end else if (bht_bank_sel_1_8_14) begin
      if (_T_10727) begin
        bht_bank_rd_data_out_1_142 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_142 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_143 <= 2'h0;
    end else if (bht_bank_sel_1_8_15) begin
      if (_T_10736) begin
        bht_bank_rd_data_out_1_143 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_143 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_144 <= 2'h0;
    end else if (bht_bank_sel_1_9_0) begin
      if (_T_10745) begin
        bht_bank_rd_data_out_1_144 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_144 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_145 <= 2'h0;
    end else if (bht_bank_sel_1_9_1) begin
      if (_T_10754) begin
        bht_bank_rd_data_out_1_145 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_145 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_146 <= 2'h0;
    end else if (bht_bank_sel_1_9_2) begin
      if (_T_10763) begin
        bht_bank_rd_data_out_1_146 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_146 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_147 <= 2'h0;
    end else if (bht_bank_sel_1_9_3) begin
      if (_T_10772) begin
        bht_bank_rd_data_out_1_147 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_147 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_148 <= 2'h0;
    end else if (bht_bank_sel_1_9_4) begin
      if (_T_10781) begin
        bht_bank_rd_data_out_1_148 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_148 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_149 <= 2'h0;
    end else if (bht_bank_sel_1_9_5) begin
      if (_T_10790) begin
        bht_bank_rd_data_out_1_149 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_149 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_150 <= 2'h0;
    end else if (bht_bank_sel_1_9_6) begin
      if (_T_10799) begin
        bht_bank_rd_data_out_1_150 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_150 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_151 <= 2'h0;
    end else if (bht_bank_sel_1_9_7) begin
      if (_T_10808) begin
        bht_bank_rd_data_out_1_151 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_151 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_152 <= 2'h0;
    end else if (bht_bank_sel_1_9_8) begin
      if (_T_10817) begin
        bht_bank_rd_data_out_1_152 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_152 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_153 <= 2'h0;
    end else if (bht_bank_sel_1_9_9) begin
      if (_T_10826) begin
        bht_bank_rd_data_out_1_153 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_153 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_154 <= 2'h0;
    end else if (bht_bank_sel_1_9_10) begin
      if (_T_10835) begin
        bht_bank_rd_data_out_1_154 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_154 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_155 <= 2'h0;
    end else if (bht_bank_sel_1_9_11) begin
      if (_T_10844) begin
        bht_bank_rd_data_out_1_155 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_155 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_156 <= 2'h0;
    end else if (bht_bank_sel_1_9_12) begin
      if (_T_10853) begin
        bht_bank_rd_data_out_1_156 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_156 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_157 <= 2'h0;
    end else if (bht_bank_sel_1_9_13) begin
      if (_T_10862) begin
        bht_bank_rd_data_out_1_157 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_157 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_158 <= 2'h0;
    end else if (bht_bank_sel_1_9_14) begin
      if (_T_10871) begin
        bht_bank_rd_data_out_1_158 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_158 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_159 <= 2'h0;
    end else if (bht_bank_sel_1_9_15) begin
      if (_T_10880) begin
        bht_bank_rd_data_out_1_159 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_159 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_160 <= 2'h0;
    end else if (bht_bank_sel_1_10_0) begin
      if (_T_10889) begin
        bht_bank_rd_data_out_1_160 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_160 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_161 <= 2'h0;
    end else if (bht_bank_sel_1_10_1) begin
      if (_T_10898) begin
        bht_bank_rd_data_out_1_161 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_161 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_162 <= 2'h0;
    end else if (bht_bank_sel_1_10_2) begin
      if (_T_10907) begin
        bht_bank_rd_data_out_1_162 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_162 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_163 <= 2'h0;
    end else if (bht_bank_sel_1_10_3) begin
      if (_T_10916) begin
        bht_bank_rd_data_out_1_163 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_163 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_164 <= 2'h0;
    end else if (bht_bank_sel_1_10_4) begin
      if (_T_10925) begin
        bht_bank_rd_data_out_1_164 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_164 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_165 <= 2'h0;
    end else if (bht_bank_sel_1_10_5) begin
      if (_T_10934) begin
        bht_bank_rd_data_out_1_165 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_165 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_166 <= 2'h0;
    end else if (bht_bank_sel_1_10_6) begin
      if (_T_10943) begin
        bht_bank_rd_data_out_1_166 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_166 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_167 <= 2'h0;
    end else if (bht_bank_sel_1_10_7) begin
      if (_T_10952) begin
        bht_bank_rd_data_out_1_167 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_167 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_168 <= 2'h0;
    end else if (bht_bank_sel_1_10_8) begin
      if (_T_10961) begin
        bht_bank_rd_data_out_1_168 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_168 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_169 <= 2'h0;
    end else if (bht_bank_sel_1_10_9) begin
      if (_T_10970) begin
        bht_bank_rd_data_out_1_169 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_169 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_170 <= 2'h0;
    end else if (bht_bank_sel_1_10_10) begin
      if (_T_10979) begin
        bht_bank_rd_data_out_1_170 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_170 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_171 <= 2'h0;
    end else if (bht_bank_sel_1_10_11) begin
      if (_T_10988) begin
        bht_bank_rd_data_out_1_171 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_171 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_172 <= 2'h0;
    end else if (bht_bank_sel_1_10_12) begin
      if (_T_10997) begin
        bht_bank_rd_data_out_1_172 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_172 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_173 <= 2'h0;
    end else if (bht_bank_sel_1_10_13) begin
      if (_T_11006) begin
        bht_bank_rd_data_out_1_173 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_173 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_174 <= 2'h0;
    end else if (bht_bank_sel_1_10_14) begin
      if (_T_11015) begin
        bht_bank_rd_data_out_1_174 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_174 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_175 <= 2'h0;
    end else if (bht_bank_sel_1_10_15) begin
      if (_T_11024) begin
        bht_bank_rd_data_out_1_175 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_175 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_176 <= 2'h0;
    end else if (bht_bank_sel_1_11_0) begin
      if (_T_11033) begin
        bht_bank_rd_data_out_1_176 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_176 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_177 <= 2'h0;
    end else if (bht_bank_sel_1_11_1) begin
      if (_T_11042) begin
        bht_bank_rd_data_out_1_177 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_177 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_178 <= 2'h0;
    end else if (bht_bank_sel_1_11_2) begin
      if (_T_11051) begin
        bht_bank_rd_data_out_1_178 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_178 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_179 <= 2'h0;
    end else if (bht_bank_sel_1_11_3) begin
      if (_T_11060) begin
        bht_bank_rd_data_out_1_179 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_179 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_180 <= 2'h0;
    end else if (bht_bank_sel_1_11_4) begin
      if (_T_11069) begin
        bht_bank_rd_data_out_1_180 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_180 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_181 <= 2'h0;
    end else if (bht_bank_sel_1_11_5) begin
      if (_T_11078) begin
        bht_bank_rd_data_out_1_181 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_181 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_182 <= 2'h0;
    end else if (bht_bank_sel_1_11_6) begin
      if (_T_11087) begin
        bht_bank_rd_data_out_1_182 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_182 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_183 <= 2'h0;
    end else if (bht_bank_sel_1_11_7) begin
      if (_T_11096) begin
        bht_bank_rd_data_out_1_183 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_183 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_184 <= 2'h0;
    end else if (bht_bank_sel_1_11_8) begin
      if (_T_11105) begin
        bht_bank_rd_data_out_1_184 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_184 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_185 <= 2'h0;
    end else if (bht_bank_sel_1_11_9) begin
      if (_T_11114) begin
        bht_bank_rd_data_out_1_185 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_185 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_186 <= 2'h0;
    end else if (bht_bank_sel_1_11_10) begin
      if (_T_11123) begin
        bht_bank_rd_data_out_1_186 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_186 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_187 <= 2'h0;
    end else if (bht_bank_sel_1_11_11) begin
      if (_T_11132) begin
        bht_bank_rd_data_out_1_187 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_187 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_188 <= 2'h0;
    end else if (bht_bank_sel_1_11_12) begin
      if (_T_11141) begin
        bht_bank_rd_data_out_1_188 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_188 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_189 <= 2'h0;
    end else if (bht_bank_sel_1_11_13) begin
      if (_T_11150) begin
        bht_bank_rd_data_out_1_189 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_189 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_190 <= 2'h0;
    end else if (bht_bank_sel_1_11_14) begin
      if (_T_11159) begin
        bht_bank_rd_data_out_1_190 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_190 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_191 <= 2'h0;
    end else if (bht_bank_sel_1_11_15) begin
      if (_T_11168) begin
        bht_bank_rd_data_out_1_191 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_191 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_192 <= 2'h0;
    end else if (bht_bank_sel_1_12_0) begin
      if (_T_11177) begin
        bht_bank_rd_data_out_1_192 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_192 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_193 <= 2'h0;
    end else if (bht_bank_sel_1_12_1) begin
      if (_T_11186) begin
        bht_bank_rd_data_out_1_193 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_193 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_194 <= 2'h0;
    end else if (bht_bank_sel_1_12_2) begin
      if (_T_11195) begin
        bht_bank_rd_data_out_1_194 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_194 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_195 <= 2'h0;
    end else if (bht_bank_sel_1_12_3) begin
      if (_T_11204) begin
        bht_bank_rd_data_out_1_195 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_195 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_196 <= 2'h0;
    end else if (bht_bank_sel_1_12_4) begin
      if (_T_11213) begin
        bht_bank_rd_data_out_1_196 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_196 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_197 <= 2'h0;
    end else if (bht_bank_sel_1_12_5) begin
      if (_T_11222) begin
        bht_bank_rd_data_out_1_197 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_197 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_198 <= 2'h0;
    end else if (bht_bank_sel_1_12_6) begin
      if (_T_11231) begin
        bht_bank_rd_data_out_1_198 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_198 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_199 <= 2'h0;
    end else if (bht_bank_sel_1_12_7) begin
      if (_T_11240) begin
        bht_bank_rd_data_out_1_199 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_199 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_200 <= 2'h0;
    end else if (bht_bank_sel_1_12_8) begin
      if (_T_11249) begin
        bht_bank_rd_data_out_1_200 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_200 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_201 <= 2'h0;
    end else if (bht_bank_sel_1_12_9) begin
      if (_T_11258) begin
        bht_bank_rd_data_out_1_201 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_201 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_202 <= 2'h0;
    end else if (bht_bank_sel_1_12_10) begin
      if (_T_11267) begin
        bht_bank_rd_data_out_1_202 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_202 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_203 <= 2'h0;
    end else if (bht_bank_sel_1_12_11) begin
      if (_T_11276) begin
        bht_bank_rd_data_out_1_203 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_203 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_204 <= 2'h0;
    end else if (bht_bank_sel_1_12_12) begin
      if (_T_11285) begin
        bht_bank_rd_data_out_1_204 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_204 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_205 <= 2'h0;
    end else if (bht_bank_sel_1_12_13) begin
      if (_T_11294) begin
        bht_bank_rd_data_out_1_205 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_205 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_206 <= 2'h0;
    end else if (bht_bank_sel_1_12_14) begin
      if (_T_11303) begin
        bht_bank_rd_data_out_1_206 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_206 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_207 <= 2'h0;
    end else if (bht_bank_sel_1_12_15) begin
      if (_T_11312) begin
        bht_bank_rd_data_out_1_207 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_207 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_208 <= 2'h0;
    end else if (bht_bank_sel_1_13_0) begin
      if (_T_11321) begin
        bht_bank_rd_data_out_1_208 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_208 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_209 <= 2'h0;
    end else if (bht_bank_sel_1_13_1) begin
      if (_T_11330) begin
        bht_bank_rd_data_out_1_209 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_209 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_210 <= 2'h0;
    end else if (bht_bank_sel_1_13_2) begin
      if (_T_11339) begin
        bht_bank_rd_data_out_1_210 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_210 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_211 <= 2'h0;
    end else if (bht_bank_sel_1_13_3) begin
      if (_T_11348) begin
        bht_bank_rd_data_out_1_211 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_211 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_212 <= 2'h0;
    end else if (bht_bank_sel_1_13_4) begin
      if (_T_11357) begin
        bht_bank_rd_data_out_1_212 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_212 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_213 <= 2'h0;
    end else if (bht_bank_sel_1_13_5) begin
      if (_T_11366) begin
        bht_bank_rd_data_out_1_213 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_213 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_214 <= 2'h0;
    end else if (bht_bank_sel_1_13_6) begin
      if (_T_11375) begin
        bht_bank_rd_data_out_1_214 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_214 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_215 <= 2'h0;
    end else if (bht_bank_sel_1_13_7) begin
      if (_T_11384) begin
        bht_bank_rd_data_out_1_215 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_215 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_216 <= 2'h0;
    end else if (bht_bank_sel_1_13_8) begin
      if (_T_11393) begin
        bht_bank_rd_data_out_1_216 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_216 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_217 <= 2'h0;
    end else if (bht_bank_sel_1_13_9) begin
      if (_T_11402) begin
        bht_bank_rd_data_out_1_217 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_217 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_218 <= 2'h0;
    end else if (bht_bank_sel_1_13_10) begin
      if (_T_11411) begin
        bht_bank_rd_data_out_1_218 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_218 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_219 <= 2'h0;
    end else if (bht_bank_sel_1_13_11) begin
      if (_T_11420) begin
        bht_bank_rd_data_out_1_219 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_219 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_220 <= 2'h0;
    end else if (bht_bank_sel_1_13_12) begin
      if (_T_11429) begin
        bht_bank_rd_data_out_1_220 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_220 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_221 <= 2'h0;
    end else if (bht_bank_sel_1_13_13) begin
      if (_T_11438) begin
        bht_bank_rd_data_out_1_221 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_221 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_222 <= 2'h0;
    end else if (bht_bank_sel_1_13_14) begin
      if (_T_11447) begin
        bht_bank_rd_data_out_1_222 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_222 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_223 <= 2'h0;
    end else if (bht_bank_sel_1_13_15) begin
      if (_T_11456) begin
        bht_bank_rd_data_out_1_223 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_223 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_224 <= 2'h0;
    end else if (bht_bank_sel_1_14_0) begin
      if (_T_11465) begin
        bht_bank_rd_data_out_1_224 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_224 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_225 <= 2'h0;
    end else if (bht_bank_sel_1_14_1) begin
      if (_T_11474) begin
        bht_bank_rd_data_out_1_225 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_225 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_226 <= 2'h0;
    end else if (bht_bank_sel_1_14_2) begin
      if (_T_11483) begin
        bht_bank_rd_data_out_1_226 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_226 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_227 <= 2'h0;
    end else if (bht_bank_sel_1_14_3) begin
      if (_T_11492) begin
        bht_bank_rd_data_out_1_227 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_227 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_228 <= 2'h0;
    end else if (bht_bank_sel_1_14_4) begin
      if (_T_11501) begin
        bht_bank_rd_data_out_1_228 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_228 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_229 <= 2'h0;
    end else if (bht_bank_sel_1_14_5) begin
      if (_T_11510) begin
        bht_bank_rd_data_out_1_229 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_229 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_230 <= 2'h0;
    end else if (bht_bank_sel_1_14_6) begin
      if (_T_11519) begin
        bht_bank_rd_data_out_1_230 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_230 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_231 <= 2'h0;
    end else if (bht_bank_sel_1_14_7) begin
      if (_T_11528) begin
        bht_bank_rd_data_out_1_231 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_231 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_232 <= 2'h0;
    end else if (bht_bank_sel_1_14_8) begin
      if (_T_11537) begin
        bht_bank_rd_data_out_1_232 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_232 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_233 <= 2'h0;
    end else if (bht_bank_sel_1_14_9) begin
      if (_T_11546) begin
        bht_bank_rd_data_out_1_233 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_233 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_234 <= 2'h0;
    end else if (bht_bank_sel_1_14_10) begin
      if (_T_11555) begin
        bht_bank_rd_data_out_1_234 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_234 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_235 <= 2'h0;
    end else if (bht_bank_sel_1_14_11) begin
      if (_T_11564) begin
        bht_bank_rd_data_out_1_235 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_235 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_236 <= 2'h0;
    end else if (bht_bank_sel_1_14_12) begin
      if (_T_11573) begin
        bht_bank_rd_data_out_1_236 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_236 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_237 <= 2'h0;
    end else if (bht_bank_sel_1_14_13) begin
      if (_T_11582) begin
        bht_bank_rd_data_out_1_237 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_237 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_238 <= 2'h0;
    end else if (bht_bank_sel_1_14_14) begin
      if (_T_11591) begin
        bht_bank_rd_data_out_1_238 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_238 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_239 <= 2'h0;
    end else if (bht_bank_sel_1_14_15) begin
      if (_T_11600) begin
        bht_bank_rd_data_out_1_239 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_239 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_240 <= 2'h0;
    end else if (bht_bank_sel_1_15_0) begin
      if (_T_11609) begin
        bht_bank_rd_data_out_1_240 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_240 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_241 <= 2'h0;
    end else if (bht_bank_sel_1_15_1) begin
      if (_T_11618) begin
        bht_bank_rd_data_out_1_241 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_241 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_242 <= 2'h0;
    end else if (bht_bank_sel_1_15_2) begin
      if (_T_11627) begin
        bht_bank_rd_data_out_1_242 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_242 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_243 <= 2'h0;
    end else if (bht_bank_sel_1_15_3) begin
      if (_T_11636) begin
        bht_bank_rd_data_out_1_243 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_243 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_244 <= 2'h0;
    end else if (bht_bank_sel_1_15_4) begin
      if (_T_11645) begin
        bht_bank_rd_data_out_1_244 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_244 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_245 <= 2'h0;
    end else if (bht_bank_sel_1_15_5) begin
      if (_T_11654) begin
        bht_bank_rd_data_out_1_245 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_245 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_246 <= 2'h0;
    end else if (bht_bank_sel_1_15_6) begin
      if (_T_11663) begin
        bht_bank_rd_data_out_1_246 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_246 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_247 <= 2'h0;
    end else if (bht_bank_sel_1_15_7) begin
      if (_T_11672) begin
        bht_bank_rd_data_out_1_247 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_247 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_248 <= 2'h0;
    end else if (bht_bank_sel_1_15_8) begin
      if (_T_11681) begin
        bht_bank_rd_data_out_1_248 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_248 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_249 <= 2'h0;
    end else if (bht_bank_sel_1_15_9) begin
      if (_T_11690) begin
        bht_bank_rd_data_out_1_249 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_249 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_250 <= 2'h0;
    end else if (bht_bank_sel_1_15_10) begin
      if (_T_11699) begin
        bht_bank_rd_data_out_1_250 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_250 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_251 <= 2'h0;
    end else if (bht_bank_sel_1_15_11) begin
      if (_T_11708) begin
        bht_bank_rd_data_out_1_251 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_251 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_252 <= 2'h0;
    end else if (bht_bank_sel_1_15_12) begin
      if (_T_11717) begin
        bht_bank_rd_data_out_1_252 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_252 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_253 <= 2'h0;
    end else if (bht_bank_sel_1_15_13) begin
      if (_T_11726) begin
        bht_bank_rd_data_out_1_253 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_253 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_254 <= 2'h0;
    end else if (bht_bank_sel_1_15_14) begin
      if (_T_11735) begin
        bht_bank_rd_data_out_1_254 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_254 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_255 <= 2'h0;
    end else if (bht_bank_sel_1_15_15) begin
      if (_T_11744) begin
        bht_bank_rd_data_out_1_255 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_255 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_0 <= 2'h0;
    end else if (bht_bank_sel_0_0_0) begin
      if (_T_7145) begin
        bht_bank_rd_data_out_0_0 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_0 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_1 <= 2'h0;
    end else if (bht_bank_sel_0_0_1) begin
      if (_T_7154) begin
        bht_bank_rd_data_out_0_1 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_1 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_2 <= 2'h0;
    end else if (bht_bank_sel_0_0_2) begin
      if (_T_7163) begin
        bht_bank_rd_data_out_0_2 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_2 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_3 <= 2'h0;
    end else if (bht_bank_sel_0_0_3) begin
      if (_T_7172) begin
        bht_bank_rd_data_out_0_3 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_3 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_4 <= 2'h0;
    end else if (bht_bank_sel_0_0_4) begin
      if (_T_7181) begin
        bht_bank_rd_data_out_0_4 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_4 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_5 <= 2'h0;
    end else if (bht_bank_sel_0_0_5) begin
      if (_T_7190) begin
        bht_bank_rd_data_out_0_5 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_5 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_6 <= 2'h0;
    end else if (bht_bank_sel_0_0_6) begin
      if (_T_7199) begin
        bht_bank_rd_data_out_0_6 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_6 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_7 <= 2'h0;
    end else if (bht_bank_sel_0_0_7) begin
      if (_T_7208) begin
        bht_bank_rd_data_out_0_7 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_7 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_8 <= 2'h0;
    end else if (bht_bank_sel_0_0_8) begin
      if (_T_7217) begin
        bht_bank_rd_data_out_0_8 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_8 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_9 <= 2'h0;
    end else if (bht_bank_sel_0_0_9) begin
      if (_T_7226) begin
        bht_bank_rd_data_out_0_9 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_9 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_10 <= 2'h0;
    end else if (bht_bank_sel_0_0_10) begin
      if (_T_7235) begin
        bht_bank_rd_data_out_0_10 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_10 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_11 <= 2'h0;
    end else if (bht_bank_sel_0_0_11) begin
      if (_T_7244) begin
        bht_bank_rd_data_out_0_11 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_11 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_12 <= 2'h0;
    end else if (bht_bank_sel_0_0_12) begin
      if (_T_7253) begin
        bht_bank_rd_data_out_0_12 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_12 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_13 <= 2'h0;
    end else if (bht_bank_sel_0_0_13) begin
      if (_T_7262) begin
        bht_bank_rd_data_out_0_13 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_13 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_14 <= 2'h0;
    end else if (bht_bank_sel_0_0_14) begin
      if (_T_7271) begin
        bht_bank_rd_data_out_0_14 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_14 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_15 <= 2'h0;
    end else if (bht_bank_sel_0_0_15) begin
      if (_T_7280) begin
        bht_bank_rd_data_out_0_15 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_15 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_16 <= 2'h0;
    end else if (bht_bank_sel_0_1_0) begin
      if (_T_7289) begin
        bht_bank_rd_data_out_0_16 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_16 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_17 <= 2'h0;
    end else if (bht_bank_sel_0_1_1) begin
      if (_T_7298) begin
        bht_bank_rd_data_out_0_17 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_17 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_18 <= 2'h0;
    end else if (bht_bank_sel_0_1_2) begin
      if (_T_7307) begin
        bht_bank_rd_data_out_0_18 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_18 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_19 <= 2'h0;
    end else if (bht_bank_sel_0_1_3) begin
      if (_T_7316) begin
        bht_bank_rd_data_out_0_19 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_19 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_20 <= 2'h0;
    end else if (bht_bank_sel_0_1_4) begin
      if (_T_7325) begin
        bht_bank_rd_data_out_0_20 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_20 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_21 <= 2'h0;
    end else if (bht_bank_sel_0_1_5) begin
      if (_T_7334) begin
        bht_bank_rd_data_out_0_21 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_21 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_22 <= 2'h0;
    end else if (bht_bank_sel_0_1_6) begin
      if (_T_7343) begin
        bht_bank_rd_data_out_0_22 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_22 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_23 <= 2'h0;
    end else if (bht_bank_sel_0_1_7) begin
      if (_T_7352) begin
        bht_bank_rd_data_out_0_23 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_23 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_24 <= 2'h0;
    end else if (bht_bank_sel_0_1_8) begin
      if (_T_7361) begin
        bht_bank_rd_data_out_0_24 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_24 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_25 <= 2'h0;
    end else if (bht_bank_sel_0_1_9) begin
      if (_T_7370) begin
        bht_bank_rd_data_out_0_25 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_25 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_26 <= 2'h0;
    end else if (bht_bank_sel_0_1_10) begin
      if (_T_7379) begin
        bht_bank_rd_data_out_0_26 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_26 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_27 <= 2'h0;
    end else if (bht_bank_sel_0_1_11) begin
      if (_T_7388) begin
        bht_bank_rd_data_out_0_27 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_27 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_28 <= 2'h0;
    end else if (bht_bank_sel_0_1_12) begin
      if (_T_7397) begin
        bht_bank_rd_data_out_0_28 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_28 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_29 <= 2'h0;
    end else if (bht_bank_sel_0_1_13) begin
      if (_T_7406) begin
        bht_bank_rd_data_out_0_29 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_29 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_30 <= 2'h0;
    end else if (bht_bank_sel_0_1_14) begin
      if (_T_7415) begin
        bht_bank_rd_data_out_0_30 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_30 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_31 <= 2'h0;
    end else if (bht_bank_sel_0_1_15) begin
      if (_T_7424) begin
        bht_bank_rd_data_out_0_31 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_31 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_32 <= 2'h0;
    end else if (bht_bank_sel_0_2_0) begin
      if (_T_7433) begin
        bht_bank_rd_data_out_0_32 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_32 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_33 <= 2'h0;
    end else if (bht_bank_sel_0_2_1) begin
      if (_T_7442) begin
        bht_bank_rd_data_out_0_33 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_33 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_34 <= 2'h0;
    end else if (bht_bank_sel_0_2_2) begin
      if (_T_7451) begin
        bht_bank_rd_data_out_0_34 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_34 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_35 <= 2'h0;
    end else if (bht_bank_sel_0_2_3) begin
      if (_T_7460) begin
        bht_bank_rd_data_out_0_35 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_35 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_36 <= 2'h0;
    end else if (bht_bank_sel_0_2_4) begin
      if (_T_7469) begin
        bht_bank_rd_data_out_0_36 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_36 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_37 <= 2'h0;
    end else if (bht_bank_sel_0_2_5) begin
      if (_T_7478) begin
        bht_bank_rd_data_out_0_37 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_37 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_38 <= 2'h0;
    end else if (bht_bank_sel_0_2_6) begin
      if (_T_7487) begin
        bht_bank_rd_data_out_0_38 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_38 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_39 <= 2'h0;
    end else if (bht_bank_sel_0_2_7) begin
      if (_T_7496) begin
        bht_bank_rd_data_out_0_39 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_39 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_40 <= 2'h0;
    end else if (bht_bank_sel_0_2_8) begin
      if (_T_7505) begin
        bht_bank_rd_data_out_0_40 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_40 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_41 <= 2'h0;
    end else if (bht_bank_sel_0_2_9) begin
      if (_T_7514) begin
        bht_bank_rd_data_out_0_41 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_41 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_42 <= 2'h0;
    end else if (bht_bank_sel_0_2_10) begin
      if (_T_7523) begin
        bht_bank_rd_data_out_0_42 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_42 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_43 <= 2'h0;
    end else if (bht_bank_sel_0_2_11) begin
      if (_T_7532) begin
        bht_bank_rd_data_out_0_43 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_43 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_44 <= 2'h0;
    end else if (bht_bank_sel_0_2_12) begin
      if (_T_7541) begin
        bht_bank_rd_data_out_0_44 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_44 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_45 <= 2'h0;
    end else if (bht_bank_sel_0_2_13) begin
      if (_T_7550) begin
        bht_bank_rd_data_out_0_45 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_45 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_46 <= 2'h0;
    end else if (bht_bank_sel_0_2_14) begin
      if (_T_7559) begin
        bht_bank_rd_data_out_0_46 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_46 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_47 <= 2'h0;
    end else if (bht_bank_sel_0_2_15) begin
      if (_T_7568) begin
        bht_bank_rd_data_out_0_47 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_47 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_48 <= 2'h0;
    end else if (bht_bank_sel_0_3_0) begin
      if (_T_7577) begin
        bht_bank_rd_data_out_0_48 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_48 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_49 <= 2'h0;
    end else if (bht_bank_sel_0_3_1) begin
      if (_T_7586) begin
        bht_bank_rd_data_out_0_49 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_49 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_50 <= 2'h0;
    end else if (bht_bank_sel_0_3_2) begin
      if (_T_7595) begin
        bht_bank_rd_data_out_0_50 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_50 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_51 <= 2'h0;
    end else if (bht_bank_sel_0_3_3) begin
      if (_T_7604) begin
        bht_bank_rd_data_out_0_51 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_51 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_52 <= 2'h0;
    end else if (bht_bank_sel_0_3_4) begin
      if (_T_7613) begin
        bht_bank_rd_data_out_0_52 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_52 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_53 <= 2'h0;
    end else if (bht_bank_sel_0_3_5) begin
      if (_T_7622) begin
        bht_bank_rd_data_out_0_53 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_53 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_54 <= 2'h0;
    end else if (bht_bank_sel_0_3_6) begin
      if (_T_7631) begin
        bht_bank_rd_data_out_0_54 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_54 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_55 <= 2'h0;
    end else if (bht_bank_sel_0_3_7) begin
      if (_T_7640) begin
        bht_bank_rd_data_out_0_55 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_55 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_56 <= 2'h0;
    end else if (bht_bank_sel_0_3_8) begin
      if (_T_7649) begin
        bht_bank_rd_data_out_0_56 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_56 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_57 <= 2'h0;
    end else if (bht_bank_sel_0_3_9) begin
      if (_T_7658) begin
        bht_bank_rd_data_out_0_57 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_57 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_58 <= 2'h0;
    end else if (bht_bank_sel_0_3_10) begin
      if (_T_7667) begin
        bht_bank_rd_data_out_0_58 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_58 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_59 <= 2'h0;
    end else if (bht_bank_sel_0_3_11) begin
      if (_T_7676) begin
        bht_bank_rd_data_out_0_59 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_59 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_60 <= 2'h0;
    end else if (bht_bank_sel_0_3_12) begin
      if (_T_7685) begin
        bht_bank_rd_data_out_0_60 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_60 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_61 <= 2'h0;
    end else if (bht_bank_sel_0_3_13) begin
      if (_T_7694) begin
        bht_bank_rd_data_out_0_61 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_61 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_62 <= 2'h0;
    end else if (bht_bank_sel_0_3_14) begin
      if (_T_7703) begin
        bht_bank_rd_data_out_0_62 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_62 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_63 <= 2'h0;
    end else if (bht_bank_sel_0_3_15) begin
      if (_T_7712) begin
        bht_bank_rd_data_out_0_63 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_63 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_64 <= 2'h0;
    end else if (bht_bank_sel_0_4_0) begin
      if (_T_7721) begin
        bht_bank_rd_data_out_0_64 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_64 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_65 <= 2'h0;
    end else if (bht_bank_sel_0_4_1) begin
      if (_T_7730) begin
        bht_bank_rd_data_out_0_65 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_65 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_66 <= 2'h0;
    end else if (bht_bank_sel_0_4_2) begin
      if (_T_7739) begin
        bht_bank_rd_data_out_0_66 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_66 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_67 <= 2'h0;
    end else if (bht_bank_sel_0_4_3) begin
      if (_T_7748) begin
        bht_bank_rd_data_out_0_67 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_67 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_68 <= 2'h0;
    end else if (bht_bank_sel_0_4_4) begin
      if (_T_7757) begin
        bht_bank_rd_data_out_0_68 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_68 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_69 <= 2'h0;
    end else if (bht_bank_sel_0_4_5) begin
      if (_T_7766) begin
        bht_bank_rd_data_out_0_69 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_69 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_70 <= 2'h0;
    end else if (bht_bank_sel_0_4_6) begin
      if (_T_7775) begin
        bht_bank_rd_data_out_0_70 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_70 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_71 <= 2'h0;
    end else if (bht_bank_sel_0_4_7) begin
      if (_T_7784) begin
        bht_bank_rd_data_out_0_71 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_71 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_72 <= 2'h0;
    end else if (bht_bank_sel_0_4_8) begin
      if (_T_7793) begin
        bht_bank_rd_data_out_0_72 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_72 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_73 <= 2'h0;
    end else if (bht_bank_sel_0_4_9) begin
      if (_T_7802) begin
        bht_bank_rd_data_out_0_73 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_73 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_74 <= 2'h0;
    end else if (bht_bank_sel_0_4_10) begin
      if (_T_7811) begin
        bht_bank_rd_data_out_0_74 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_74 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_75 <= 2'h0;
    end else if (bht_bank_sel_0_4_11) begin
      if (_T_7820) begin
        bht_bank_rd_data_out_0_75 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_75 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_76 <= 2'h0;
    end else if (bht_bank_sel_0_4_12) begin
      if (_T_7829) begin
        bht_bank_rd_data_out_0_76 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_76 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_77 <= 2'h0;
    end else if (bht_bank_sel_0_4_13) begin
      if (_T_7838) begin
        bht_bank_rd_data_out_0_77 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_77 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_78 <= 2'h0;
    end else if (bht_bank_sel_0_4_14) begin
      if (_T_7847) begin
        bht_bank_rd_data_out_0_78 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_78 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_79 <= 2'h0;
    end else if (bht_bank_sel_0_4_15) begin
      if (_T_7856) begin
        bht_bank_rd_data_out_0_79 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_79 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_80 <= 2'h0;
    end else if (bht_bank_sel_0_5_0) begin
      if (_T_7865) begin
        bht_bank_rd_data_out_0_80 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_80 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_81 <= 2'h0;
    end else if (bht_bank_sel_0_5_1) begin
      if (_T_7874) begin
        bht_bank_rd_data_out_0_81 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_81 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_82 <= 2'h0;
    end else if (bht_bank_sel_0_5_2) begin
      if (_T_7883) begin
        bht_bank_rd_data_out_0_82 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_82 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_83 <= 2'h0;
    end else if (bht_bank_sel_0_5_3) begin
      if (_T_7892) begin
        bht_bank_rd_data_out_0_83 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_83 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_84 <= 2'h0;
    end else if (bht_bank_sel_0_5_4) begin
      if (_T_7901) begin
        bht_bank_rd_data_out_0_84 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_84 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_85 <= 2'h0;
    end else if (bht_bank_sel_0_5_5) begin
      if (_T_7910) begin
        bht_bank_rd_data_out_0_85 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_85 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_86 <= 2'h0;
    end else if (bht_bank_sel_0_5_6) begin
      if (_T_7919) begin
        bht_bank_rd_data_out_0_86 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_86 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_87 <= 2'h0;
    end else if (bht_bank_sel_0_5_7) begin
      if (_T_7928) begin
        bht_bank_rd_data_out_0_87 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_87 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_88 <= 2'h0;
    end else if (bht_bank_sel_0_5_8) begin
      if (_T_7937) begin
        bht_bank_rd_data_out_0_88 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_88 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_89 <= 2'h0;
    end else if (bht_bank_sel_0_5_9) begin
      if (_T_7946) begin
        bht_bank_rd_data_out_0_89 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_89 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_90 <= 2'h0;
    end else if (bht_bank_sel_0_5_10) begin
      if (_T_7955) begin
        bht_bank_rd_data_out_0_90 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_90 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_91 <= 2'h0;
    end else if (bht_bank_sel_0_5_11) begin
      if (_T_7964) begin
        bht_bank_rd_data_out_0_91 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_91 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_92 <= 2'h0;
    end else if (bht_bank_sel_0_5_12) begin
      if (_T_7973) begin
        bht_bank_rd_data_out_0_92 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_92 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_93 <= 2'h0;
    end else if (bht_bank_sel_0_5_13) begin
      if (_T_7982) begin
        bht_bank_rd_data_out_0_93 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_93 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_94 <= 2'h0;
    end else if (bht_bank_sel_0_5_14) begin
      if (_T_7991) begin
        bht_bank_rd_data_out_0_94 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_94 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_95 <= 2'h0;
    end else if (bht_bank_sel_0_5_15) begin
      if (_T_8000) begin
        bht_bank_rd_data_out_0_95 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_95 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_96 <= 2'h0;
    end else if (bht_bank_sel_0_6_0) begin
      if (_T_8009) begin
        bht_bank_rd_data_out_0_96 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_96 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_97 <= 2'h0;
    end else if (bht_bank_sel_0_6_1) begin
      if (_T_8018) begin
        bht_bank_rd_data_out_0_97 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_97 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_98 <= 2'h0;
    end else if (bht_bank_sel_0_6_2) begin
      if (_T_8027) begin
        bht_bank_rd_data_out_0_98 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_98 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_99 <= 2'h0;
    end else if (bht_bank_sel_0_6_3) begin
      if (_T_8036) begin
        bht_bank_rd_data_out_0_99 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_99 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_100 <= 2'h0;
    end else if (bht_bank_sel_0_6_4) begin
      if (_T_8045) begin
        bht_bank_rd_data_out_0_100 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_100 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_101 <= 2'h0;
    end else if (bht_bank_sel_0_6_5) begin
      if (_T_8054) begin
        bht_bank_rd_data_out_0_101 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_101 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_102 <= 2'h0;
    end else if (bht_bank_sel_0_6_6) begin
      if (_T_8063) begin
        bht_bank_rd_data_out_0_102 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_102 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_103 <= 2'h0;
    end else if (bht_bank_sel_0_6_7) begin
      if (_T_8072) begin
        bht_bank_rd_data_out_0_103 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_103 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_104 <= 2'h0;
    end else if (bht_bank_sel_0_6_8) begin
      if (_T_8081) begin
        bht_bank_rd_data_out_0_104 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_104 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_105 <= 2'h0;
    end else if (bht_bank_sel_0_6_9) begin
      if (_T_8090) begin
        bht_bank_rd_data_out_0_105 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_105 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_106 <= 2'h0;
    end else if (bht_bank_sel_0_6_10) begin
      if (_T_8099) begin
        bht_bank_rd_data_out_0_106 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_106 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_107 <= 2'h0;
    end else if (bht_bank_sel_0_6_11) begin
      if (_T_8108) begin
        bht_bank_rd_data_out_0_107 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_107 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_108 <= 2'h0;
    end else if (bht_bank_sel_0_6_12) begin
      if (_T_8117) begin
        bht_bank_rd_data_out_0_108 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_108 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_109 <= 2'h0;
    end else if (bht_bank_sel_0_6_13) begin
      if (_T_8126) begin
        bht_bank_rd_data_out_0_109 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_109 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_110 <= 2'h0;
    end else if (bht_bank_sel_0_6_14) begin
      if (_T_8135) begin
        bht_bank_rd_data_out_0_110 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_110 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_111 <= 2'h0;
    end else if (bht_bank_sel_0_6_15) begin
      if (_T_8144) begin
        bht_bank_rd_data_out_0_111 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_111 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_112 <= 2'h0;
    end else if (bht_bank_sel_0_7_0) begin
      if (_T_8153) begin
        bht_bank_rd_data_out_0_112 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_112 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_113 <= 2'h0;
    end else if (bht_bank_sel_0_7_1) begin
      if (_T_8162) begin
        bht_bank_rd_data_out_0_113 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_113 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_114 <= 2'h0;
    end else if (bht_bank_sel_0_7_2) begin
      if (_T_8171) begin
        bht_bank_rd_data_out_0_114 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_114 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_115 <= 2'h0;
    end else if (bht_bank_sel_0_7_3) begin
      if (_T_8180) begin
        bht_bank_rd_data_out_0_115 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_115 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_116 <= 2'h0;
    end else if (bht_bank_sel_0_7_4) begin
      if (_T_8189) begin
        bht_bank_rd_data_out_0_116 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_116 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_117 <= 2'h0;
    end else if (bht_bank_sel_0_7_5) begin
      if (_T_8198) begin
        bht_bank_rd_data_out_0_117 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_117 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_118 <= 2'h0;
    end else if (bht_bank_sel_0_7_6) begin
      if (_T_8207) begin
        bht_bank_rd_data_out_0_118 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_118 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_119 <= 2'h0;
    end else if (bht_bank_sel_0_7_7) begin
      if (_T_8216) begin
        bht_bank_rd_data_out_0_119 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_119 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_120 <= 2'h0;
    end else if (bht_bank_sel_0_7_8) begin
      if (_T_8225) begin
        bht_bank_rd_data_out_0_120 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_120 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_121 <= 2'h0;
    end else if (bht_bank_sel_0_7_9) begin
      if (_T_8234) begin
        bht_bank_rd_data_out_0_121 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_121 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_122 <= 2'h0;
    end else if (bht_bank_sel_0_7_10) begin
      if (_T_8243) begin
        bht_bank_rd_data_out_0_122 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_122 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_123 <= 2'h0;
    end else if (bht_bank_sel_0_7_11) begin
      if (_T_8252) begin
        bht_bank_rd_data_out_0_123 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_123 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_124 <= 2'h0;
    end else if (bht_bank_sel_0_7_12) begin
      if (_T_8261) begin
        bht_bank_rd_data_out_0_124 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_124 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_125 <= 2'h0;
    end else if (bht_bank_sel_0_7_13) begin
      if (_T_8270) begin
        bht_bank_rd_data_out_0_125 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_125 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_126 <= 2'h0;
    end else if (bht_bank_sel_0_7_14) begin
      if (_T_8279) begin
        bht_bank_rd_data_out_0_126 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_126 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_127 <= 2'h0;
    end else if (bht_bank_sel_0_7_15) begin
      if (_T_8288) begin
        bht_bank_rd_data_out_0_127 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_127 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_128 <= 2'h0;
    end else if (bht_bank_sel_0_8_0) begin
      if (_T_8297) begin
        bht_bank_rd_data_out_0_128 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_128 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_129 <= 2'h0;
    end else if (bht_bank_sel_0_8_1) begin
      if (_T_8306) begin
        bht_bank_rd_data_out_0_129 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_129 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_130 <= 2'h0;
    end else if (bht_bank_sel_0_8_2) begin
      if (_T_8315) begin
        bht_bank_rd_data_out_0_130 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_130 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_131 <= 2'h0;
    end else if (bht_bank_sel_0_8_3) begin
      if (_T_8324) begin
        bht_bank_rd_data_out_0_131 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_131 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_132 <= 2'h0;
    end else if (bht_bank_sel_0_8_4) begin
      if (_T_8333) begin
        bht_bank_rd_data_out_0_132 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_132 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_133 <= 2'h0;
    end else if (bht_bank_sel_0_8_5) begin
      if (_T_8342) begin
        bht_bank_rd_data_out_0_133 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_133 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_134 <= 2'h0;
    end else if (bht_bank_sel_0_8_6) begin
      if (_T_8351) begin
        bht_bank_rd_data_out_0_134 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_134 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_135 <= 2'h0;
    end else if (bht_bank_sel_0_8_7) begin
      if (_T_8360) begin
        bht_bank_rd_data_out_0_135 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_135 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_136 <= 2'h0;
    end else if (bht_bank_sel_0_8_8) begin
      if (_T_8369) begin
        bht_bank_rd_data_out_0_136 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_136 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_137 <= 2'h0;
    end else if (bht_bank_sel_0_8_9) begin
      if (_T_8378) begin
        bht_bank_rd_data_out_0_137 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_137 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_138 <= 2'h0;
    end else if (bht_bank_sel_0_8_10) begin
      if (_T_8387) begin
        bht_bank_rd_data_out_0_138 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_138 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_139 <= 2'h0;
    end else if (bht_bank_sel_0_8_11) begin
      if (_T_8396) begin
        bht_bank_rd_data_out_0_139 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_139 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_140 <= 2'h0;
    end else if (bht_bank_sel_0_8_12) begin
      if (_T_8405) begin
        bht_bank_rd_data_out_0_140 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_140 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_141 <= 2'h0;
    end else if (bht_bank_sel_0_8_13) begin
      if (_T_8414) begin
        bht_bank_rd_data_out_0_141 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_141 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_142 <= 2'h0;
    end else if (bht_bank_sel_0_8_14) begin
      if (_T_8423) begin
        bht_bank_rd_data_out_0_142 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_142 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_143 <= 2'h0;
    end else if (bht_bank_sel_0_8_15) begin
      if (_T_8432) begin
        bht_bank_rd_data_out_0_143 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_143 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_144 <= 2'h0;
    end else if (bht_bank_sel_0_9_0) begin
      if (_T_8441) begin
        bht_bank_rd_data_out_0_144 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_144 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_145 <= 2'h0;
    end else if (bht_bank_sel_0_9_1) begin
      if (_T_8450) begin
        bht_bank_rd_data_out_0_145 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_145 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_146 <= 2'h0;
    end else if (bht_bank_sel_0_9_2) begin
      if (_T_8459) begin
        bht_bank_rd_data_out_0_146 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_146 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_147 <= 2'h0;
    end else if (bht_bank_sel_0_9_3) begin
      if (_T_8468) begin
        bht_bank_rd_data_out_0_147 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_147 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_148 <= 2'h0;
    end else if (bht_bank_sel_0_9_4) begin
      if (_T_8477) begin
        bht_bank_rd_data_out_0_148 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_148 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_149 <= 2'h0;
    end else if (bht_bank_sel_0_9_5) begin
      if (_T_8486) begin
        bht_bank_rd_data_out_0_149 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_149 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_150 <= 2'h0;
    end else if (bht_bank_sel_0_9_6) begin
      if (_T_8495) begin
        bht_bank_rd_data_out_0_150 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_150 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_151 <= 2'h0;
    end else if (bht_bank_sel_0_9_7) begin
      if (_T_8504) begin
        bht_bank_rd_data_out_0_151 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_151 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_152 <= 2'h0;
    end else if (bht_bank_sel_0_9_8) begin
      if (_T_8513) begin
        bht_bank_rd_data_out_0_152 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_152 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_153 <= 2'h0;
    end else if (bht_bank_sel_0_9_9) begin
      if (_T_8522) begin
        bht_bank_rd_data_out_0_153 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_153 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_154 <= 2'h0;
    end else if (bht_bank_sel_0_9_10) begin
      if (_T_8531) begin
        bht_bank_rd_data_out_0_154 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_154 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_155 <= 2'h0;
    end else if (bht_bank_sel_0_9_11) begin
      if (_T_8540) begin
        bht_bank_rd_data_out_0_155 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_155 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_156 <= 2'h0;
    end else if (bht_bank_sel_0_9_12) begin
      if (_T_8549) begin
        bht_bank_rd_data_out_0_156 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_156 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_157 <= 2'h0;
    end else if (bht_bank_sel_0_9_13) begin
      if (_T_8558) begin
        bht_bank_rd_data_out_0_157 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_157 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_158 <= 2'h0;
    end else if (bht_bank_sel_0_9_14) begin
      if (_T_8567) begin
        bht_bank_rd_data_out_0_158 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_158 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_159 <= 2'h0;
    end else if (bht_bank_sel_0_9_15) begin
      if (_T_8576) begin
        bht_bank_rd_data_out_0_159 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_159 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_160 <= 2'h0;
    end else if (bht_bank_sel_0_10_0) begin
      if (_T_8585) begin
        bht_bank_rd_data_out_0_160 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_160 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_161 <= 2'h0;
    end else if (bht_bank_sel_0_10_1) begin
      if (_T_8594) begin
        bht_bank_rd_data_out_0_161 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_161 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_162 <= 2'h0;
    end else if (bht_bank_sel_0_10_2) begin
      if (_T_8603) begin
        bht_bank_rd_data_out_0_162 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_162 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_163 <= 2'h0;
    end else if (bht_bank_sel_0_10_3) begin
      if (_T_8612) begin
        bht_bank_rd_data_out_0_163 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_163 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_164 <= 2'h0;
    end else if (bht_bank_sel_0_10_4) begin
      if (_T_8621) begin
        bht_bank_rd_data_out_0_164 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_164 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_165 <= 2'h0;
    end else if (bht_bank_sel_0_10_5) begin
      if (_T_8630) begin
        bht_bank_rd_data_out_0_165 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_165 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_166 <= 2'h0;
    end else if (bht_bank_sel_0_10_6) begin
      if (_T_8639) begin
        bht_bank_rd_data_out_0_166 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_166 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_167 <= 2'h0;
    end else if (bht_bank_sel_0_10_7) begin
      if (_T_8648) begin
        bht_bank_rd_data_out_0_167 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_167 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_168 <= 2'h0;
    end else if (bht_bank_sel_0_10_8) begin
      if (_T_8657) begin
        bht_bank_rd_data_out_0_168 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_168 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_169 <= 2'h0;
    end else if (bht_bank_sel_0_10_9) begin
      if (_T_8666) begin
        bht_bank_rd_data_out_0_169 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_169 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_170 <= 2'h0;
    end else if (bht_bank_sel_0_10_10) begin
      if (_T_8675) begin
        bht_bank_rd_data_out_0_170 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_170 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_171 <= 2'h0;
    end else if (bht_bank_sel_0_10_11) begin
      if (_T_8684) begin
        bht_bank_rd_data_out_0_171 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_171 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_172 <= 2'h0;
    end else if (bht_bank_sel_0_10_12) begin
      if (_T_8693) begin
        bht_bank_rd_data_out_0_172 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_172 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_173 <= 2'h0;
    end else if (bht_bank_sel_0_10_13) begin
      if (_T_8702) begin
        bht_bank_rd_data_out_0_173 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_173 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_174 <= 2'h0;
    end else if (bht_bank_sel_0_10_14) begin
      if (_T_8711) begin
        bht_bank_rd_data_out_0_174 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_174 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_175 <= 2'h0;
    end else if (bht_bank_sel_0_10_15) begin
      if (_T_8720) begin
        bht_bank_rd_data_out_0_175 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_175 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_176 <= 2'h0;
    end else if (bht_bank_sel_0_11_0) begin
      if (_T_8729) begin
        bht_bank_rd_data_out_0_176 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_176 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_177 <= 2'h0;
    end else if (bht_bank_sel_0_11_1) begin
      if (_T_8738) begin
        bht_bank_rd_data_out_0_177 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_177 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_178 <= 2'h0;
    end else if (bht_bank_sel_0_11_2) begin
      if (_T_8747) begin
        bht_bank_rd_data_out_0_178 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_178 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_179 <= 2'h0;
    end else if (bht_bank_sel_0_11_3) begin
      if (_T_8756) begin
        bht_bank_rd_data_out_0_179 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_179 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_180 <= 2'h0;
    end else if (bht_bank_sel_0_11_4) begin
      if (_T_8765) begin
        bht_bank_rd_data_out_0_180 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_180 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_181 <= 2'h0;
    end else if (bht_bank_sel_0_11_5) begin
      if (_T_8774) begin
        bht_bank_rd_data_out_0_181 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_181 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_182 <= 2'h0;
    end else if (bht_bank_sel_0_11_6) begin
      if (_T_8783) begin
        bht_bank_rd_data_out_0_182 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_182 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_183 <= 2'h0;
    end else if (bht_bank_sel_0_11_7) begin
      if (_T_8792) begin
        bht_bank_rd_data_out_0_183 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_183 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_184 <= 2'h0;
    end else if (bht_bank_sel_0_11_8) begin
      if (_T_8801) begin
        bht_bank_rd_data_out_0_184 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_184 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_185 <= 2'h0;
    end else if (bht_bank_sel_0_11_9) begin
      if (_T_8810) begin
        bht_bank_rd_data_out_0_185 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_185 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_186 <= 2'h0;
    end else if (bht_bank_sel_0_11_10) begin
      if (_T_8819) begin
        bht_bank_rd_data_out_0_186 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_186 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_187 <= 2'h0;
    end else if (bht_bank_sel_0_11_11) begin
      if (_T_8828) begin
        bht_bank_rd_data_out_0_187 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_187 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_188 <= 2'h0;
    end else if (bht_bank_sel_0_11_12) begin
      if (_T_8837) begin
        bht_bank_rd_data_out_0_188 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_188 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_189 <= 2'h0;
    end else if (bht_bank_sel_0_11_13) begin
      if (_T_8846) begin
        bht_bank_rd_data_out_0_189 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_189 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_190 <= 2'h0;
    end else if (bht_bank_sel_0_11_14) begin
      if (_T_8855) begin
        bht_bank_rd_data_out_0_190 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_190 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_191 <= 2'h0;
    end else if (bht_bank_sel_0_11_15) begin
      if (_T_8864) begin
        bht_bank_rd_data_out_0_191 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_191 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_192 <= 2'h0;
    end else if (bht_bank_sel_0_12_0) begin
      if (_T_8873) begin
        bht_bank_rd_data_out_0_192 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_192 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_193 <= 2'h0;
    end else if (bht_bank_sel_0_12_1) begin
      if (_T_8882) begin
        bht_bank_rd_data_out_0_193 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_193 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_194 <= 2'h0;
    end else if (bht_bank_sel_0_12_2) begin
      if (_T_8891) begin
        bht_bank_rd_data_out_0_194 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_194 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_195 <= 2'h0;
    end else if (bht_bank_sel_0_12_3) begin
      if (_T_8900) begin
        bht_bank_rd_data_out_0_195 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_195 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_196 <= 2'h0;
    end else if (bht_bank_sel_0_12_4) begin
      if (_T_8909) begin
        bht_bank_rd_data_out_0_196 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_196 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_197 <= 2'h0;
    end else if (bht_bank_sel_0_12_5) begin
      if (_T_8918) begin
        bht_bank_rd_data_out_0_197 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_197 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_198 <= 2'h0;
    end else if (bht_bank_sel_0_12_6) begin
      if (_T_8927) begin
        bht_bank_rd_data_out_0_198 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_198 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_199 <= 2'h0;
    end else if (bht_bank_sel_0_12_7) begin
      if (_T_8936) begin
        bht_bank_rd_data_out_0_199 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_199 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_200 <= 2'h0;
    end else if (bht_bank_sel_0_12_8) begin
      if (_T_8945) begin
        bht_bank_rd_data_out_0_200 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_200 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_201 <= 2'h0;
    end else if (bht_bank_sel_0_12_9) begin
      if (_T_8954) begin
        bht_bank_rd_data_out_0_201 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_201 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_202 <= 2'h0;
    end else if (bht_bank_sel_0_12_10) begin
      if (_T_8963) begin
        bht_bank_rd_data_out_0_202 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_202 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_203 <= 2'h0;
    end else if (bht_bank_sel_0_12_11) begin
      if (_T_8972) begin
        bht_bank_rd_data_out_0_203 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_203 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_204 <= 2'h0;
    end else if (bht_bank_sel_0_12_12) begin
      if (_T_8981) begin
        bht_bank_rd_data_out_0_204 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_204 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_205 <= 2'h0;
    end else if (bht_bank_sel_0_12_13) begin
      if (_T_8990) begin
        bht_bank_rd_data_out_0_205 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_205 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_206 <= 2'h0;
    end else if (bht_bank_sel_0_12_14) begin
      if (_T_8999) begin
        bht_bank_rd_data_out_0_206 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_206 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_207 <= 2'h0;
    end else if (bht_bank_sel_0_12_15) begin
      if (_T_9008) begin
        bht_bank_rd_data_out_0_207 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_207 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_208 <= 2'h0;
    end else if (bht_bank_sel_0_13_0) begin
      if (_T_9017) begin
        bht_bank_rd_data_out_0_208 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_208 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_209 <= 2'h0;
    end else if (bht_bank_sel_0_13_1) begin
      if (_T_9026) begin
        bht_bank_rd_data_out_0_209 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_209 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_210 <= 2'h0;
    end else if (bht_bank_sel_0_13_2) begin
      if (_T_9035) begin
        bht_bank_rd_data_out_0_210 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_210 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_211 <= 2'h0;
    end else if (bht_bank_sel_0_13_3) begin
      if (_T_9044) begin
        bht_bank_rd_data_out_0_211 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_211 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_212 <= 2'h0;
    end else if (bht_bank_sel_0_13_4) begin
      if (_T_9053) begin
        bht_bank_rd_data_out_0_212 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_212 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_213 <= 2'h0;
    end else if (bht_bank_sel_0_13_5) begin
      if (_T_9062) begin
        bht_bank_rd_data_out_0_213 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_213 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_214 <= 2'h0;
    end else if (bht_bank_sel_0_13_6) begin
      if (_T_9071) begin
        bht_bank_rd_data_out_0_214 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_214 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_215 <= 2'h0;
    end else if (bht_bank_sel_0_13_7) begin
      if (_T_9080) begin
        bht_bank_rd_data_out_0_215 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_215 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_216 <= 2'h0;
    end else if (bht_bank_sel_0_13_8) begin
      if (_T_9089) begin
        bht_bank_rd_data_out_0_216 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_216 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_217 <= 2'h0;
    end else if (bht_bank_sel_0_13_9) begin
      if (_T_9098) begin
        bht_bank_rd_data_out_0_217 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_217 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_218 <= 2'h0;
    end else if (bht_bank_sel_0_13_10) begin
      if (_T_9107) begin
        bht_bank_rd_data_out_0_218 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_218 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_219 <= 2'h0;
    end else if (bht_bank_sel_0_13_11) begin
      if (_T_9116) begin
        bht_bank_rd_data_out_0_219 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_219 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_220 <= 2'h0;
    end else if (bht_bank_sel_0_13_12) begin
      if (_T_9125) begin
        bht_bank_rd_data_out_0_220 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_220 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_221 <= 2'h0;
    end else if (bht_bank_sel_0_13_13) begin
      if (_T_9134) begin
        bht_bank_rd_data_out_0_221 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_221 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_222 <= 2'h0;
    end else if (bht_bank_sel_0_13_14) begin
      if (_T_9143) begin
        bht_bank_rd_data_out_0_222 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_222 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_223 <= 2'h0;
    end else if (bht_bank_sel_0_13_15) begin
      if (_T_9152) begin
        bht_bank_rd_data_out_0_223 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_223 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_224 <= 2'h0;
    end else if (bht_bank_sel_0_14_0) begin
      if (_T_9161) begin
        bht_bank_rd_data_out_0_224 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_224 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_225 <= 2'h0;
    end else if (bht_bank_sel_0_14_1) begin
      if (_T_9170) begin
        bht_bank_rd_data_out_0_225 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_225 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_226 <= 2'h0;
    end else if (bht_bank_sel_0_14_2) begin
      if (_T_9179) begin
        bht_bank_rd_data_out_0_226 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_226 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_227 <= 2'h0;
    end else if (bht_bank_sel_0_14_3) begin
      if (_T_9188) begin
        bht_bank_rd_data_out_0_227 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_227 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_228 <= 2'h0;
    end else if (bht_bank_sel_0_14_4) begin
      if (_T_9197) begin
        bht_bank_rd_data_out_0_228 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_228 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_229 <= 2'h0;
    end else if (bht_bank_sel_0_14_5) begin
      if (_T_9206) begin
        bht_bank_rd_data_out_0_229 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_229 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_230 <= 2'h0;
    end else if (bht_bank_sel_0_14_6) begin
      if (_T_9215) begin
        bht_bank_rd_data_out_0_230 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_230 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_231 <= 2'h0;
    end else if (bht_bank_sel_0_14_7) begin
      if (_T_9224) begin
        bht_bank_rd_data_out_0_231 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_231 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_232 <= 2'h0;
    end else if (bht_bank_sel_0_14_8) begin
      if (_T_9233) begin
        bht_bank_rd_data_out_0_232 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_232 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_233 <= 2'h0;
    end else if (bht_bank_sel_0_14_9) begin
      if (_T_9242) begin
        bht_bank_rd_data_out_0_233 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_233 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_234 <= 2'h0;
    end else if (bht_bank_sel_0_14_10) begin
      if (_T_9251) begin
        bht_bank_rd_data_out_0_234 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_234 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_235 <= 2'h0;
    end else if (bht_bank_sel_0_14_11) begin
      if (_T_9260) begin
        bht_bank_rd_data_out_0_235 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_235 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_236 <= 2'h0;
    end else if (bht_bank_sel_0_14_12) begin
      if (_T_9269) begin
        bht_bank_rd_data_out_0_236 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_236 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_237 <= 2'h0;
    end else if (bht_bank_sel_0_14_13) begin
      if (_T_9278) begin
        bht_bank_rd_data_out_0_237 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_237 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_238 <= 2'h0;
    end else if (bht_bank_sel_0_14_14) begin
      if (_T_9287) begin
        bht_bank_rd_data_out_0_238 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_238 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_239 <= 2'h0;
    end else if (bht_bank_sel_0_14_15) begin
      if (_T_9296) begin
        bht_bank_rd_data_out_0_239 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_239 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_240 <= 2'h0;
    end else if (bht_bank_sel_0_15_0) begin
      if (_T_9305) begin
        bht_bank_rd_data_out_0_240 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_240 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_241 <= 2'h0;
    end else if (bht_bank_sel_0_15_1) begin
      if (_T_9314) begin
        bht_bank_rd_data_out_0_241 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_241 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_242 <= 2'h0;
    end else if (bht_bank_sel_0_15_2) begin
      if (_T_9323) begin
        bht_bank_rd_data_out_0_242 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_242 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_243 <= 2'h0;
    end else if (bht_bank_sel_0_15_3) begin
      if (_T_9332) begin
        bht_bank_rd_data_out_0_243 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_243 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_244 <= 2'h0;
    end else if (bht_bank_sel_0_15_4) begin
      if (_T_9341) begin
        bht_bank_rd_data_out_0_244 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_244 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_245 <= 2'h0;
    end else if (bht_bank_sel_0_15_5) begin
      if (_T_9350) begin
        bht_bank_rd_data_out_0_245 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_245 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_246 <= 2'h0;
    end else if (bht_bank_sel_0_15_6) begin
      if (_T_9359) begin
        bht_bank_rd_data_out_0_246 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_246 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_247 <= 2'h0;
    end else if (bht_bank_sel_0_15_7) begin
      if (_T_9368) begin
        bht_bank_rd_data_out_0_247 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_247 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_248 <= 2'h0;
    end else if (bht_bank_sel_0_15_8) begin
      if (_T_9377) begin
        bht_bank_rd_data_out_0_248 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_248 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_249 <= 2'h0;
    end else if (bht_bank_sel_0_15_9) begin
      if (_T_9386) begin
        bht_bank_rd_data_out_0_249 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_249 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_250 <= 2'h0;
    end else if (bht_bank_sel_0_15_10) begin
      if (_T_9395) begin
        bht_bank_rd_data_out_0_250 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_250 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_251 <= 2'h0;
    end else if (bht_bank_sel_0_15_11) begin
      if (_T_9404) begin
        bht_bank_rd_data_out_0_251 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_251 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_252 <= 2'h0;
    end else if (bht_bank_sel_0_15_12) begin
      if (_T_9413) begin
        bht_bank_rd_data_out_0_252 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_252 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_253 <= 2'h0;
    end else if (bht_bank_sel_0_15_13) begin
      if (_T_9422) begin
        bht_bank_rd_data_out_0_253 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_253 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_254 <= 2'h0;
    end else if (bht_bank_sel_0_15_14) begin
      if (_T_9431) begin
        bht_bank_rd_data_out_0_254 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_254 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_255 <= 2'h0;
    end else if (bht_bank_sel_0_15_15) begin
      if (_T_9440) begin
        bht_bank_rd_data_out_0_255 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_255 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      exu_mp_way_f <= 1'h0;
    end else if (_T_367) begin
      exu_mp_way_f <= io_exu_bp_exu_mp_pkt_bits_way;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_lru_b0_f <= 256'h0;
    end else if (_T_234) begin
      btb_lru_b0_f <= _T_203;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      exu_flush_final_d1 <= 1'h0;
    end else if (_T_371) begin
      exu_flush_final_d1 <= io_exu_flush_final;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifc_fetch_adder_prior <= 30'h0;
    end else if (_T_411) begin
      ifc_fetch_adder_prior <= io_ifc_fetch_addr_f[30:1];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_0 <= 32'h0;
    end else if (rsenable_0) begin
      rets_out_0 <= rets_in_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_1 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_1 <= rets_in_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_2 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_2 <= rets_in_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_3 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_3 <= rets_in_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_4 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_4 <= rets_in_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_5 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_5 <= rets_in_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_6 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_6 <= rets_in_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_7 <= 32'h0;
    end else if (rs_push) begin
      rets_out_7 <= rets_out_6;
    end
  end
endmodule
module ifu_compress_ctl(
  input  [15:0] io_din,
  output [31:0] io_dout
);
  wire  _T_2 = ~io_din[14]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_4 = ~io_din[13]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_7 = ~io_din[6]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_9 = ~io_din[5]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_11 = io_din[15] & _T_2; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_12 = _T_11 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_13 = _T_12 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_14 = _T_13 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_15 = _T_14 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_16 = _T_15 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_23 = ~io_din[11]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_28 = _T_12 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_29 = _T_28 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_30 = _T_29 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_30 = _T_16 | _T_30; // @[ifu_compress_ctl.scala 17:53]
  wire  _T_38 = ~io_din[10]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_40 = ~io_din[9]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_42 = ~io_din[8]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_44 = ~io_din[7]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_50 = ~io_din[4]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_52 = ~io_din[3]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_54 = ~io_din[2]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_56 = _T_2 & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_57 = _T_56 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_58 = _T_57 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_59 = _T_58 & _T_40; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_60 = _T_59 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_61 = _T_60 & _T_44; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_62 = _T_61 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_63 = _T_62 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_64 = _T_63 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_65 = _T_64 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_66 = _T_65 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  out_20 = _T_66 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_79 = _T_28 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_90 = _T_12 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_91 = _T_90 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_92 = _T_79 | _T_91; // @[ifu_compress_ctl.scala 21:46]
  wire  _T_102 = _T_12 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_103 = _T_102 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_104 = _T_92 | _T_103; // @[ifu_compress_ctl.scala 21:80]
  wire  _T_114 = _T_12 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_115 = _T_114 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_14 = _T_104 | _T_115; // @[ifu_compress_ctl.scala 21:113]
  wire  _T_128 = _T_12 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_129 = _T_128 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_130 = _T_129 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_142 = _T_128 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_143 = _T_142 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_144 = _T_130 | _T_143; // @[ifu_compress_ctl.scala 23:50]
  wire  _T_147 = ~io_din[0]; // @[ifu_compress_ctl.scala 23:101]
  wire  _T_148 = io_din[14] & _T_147; // @[ifu_compress_ctl.scala 23:99]
  wire  out_13 = _T_144 | _T_148; // @[ifu_compress_ctl.scala 23:86]
  wire  _T_161 = _T_102 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_162 = _T_161 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_175 = _T_162 | _T_79; // @[ifu_compress_ctl.scala 25:47]
  wire  _T_188 = _T_175 | _T_91; // @[ifu_compress_ctl.scala 25:81]
  wire  _T_190 = ~io_din[15]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_194 = _T_190 & _T_2; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_195 = _T_194 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_196 = _T_188 | _T_195; // @[ifu_compress_ctl.scala 25:115]
  wire  _T_200 = io_din[15] & io_din[14]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_201 = _T_200 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_12 = _T_196 | _T_201; // @[ifu_compress_ctl.scala 26:26]
  wire  _T_217 = _T_11 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_218 = _T_217 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_219 = _T_218 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_220 = _T_219 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_221 = _T_220 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_224 = _T_221 & _T_147; // @[ifu_compress_ctl.scala 28:53]
  wire  _T_228 = _T_2 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_229 = _T_224 | _T_228; // @[ifu_compress_ctl.scala 28:67]
  wire  _T_234 = _T_200 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_6 = _T_229 | _T_234; // @[ifu_compress_ctl.scala 28:88]
  wire  _T_239 = io_din[15] & _T_147; // @[ifu_compress_ctl.scala 30:24]
  wire  _T_243 = io_din[15] & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_244 = _T_243 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_245 = _T_239 | _T_244; // @[ifu_compress_ctl.scala 30:39]
  wire  _T_249 = io_din[13] & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_250 = _T_245 | _T_249; // @[ifu_compress_ctl.scala 30:63]
  wire  _T_253 = io_din[13] & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_254 = _T_250 | _T_253; // @[ifu_compress_ctl.scala 30:83]
  wire  _T_257 = io_din[13] & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_258 = _T_254 | _T_257; // @[ifu_compress_ctl.scala 30:102]
  wire  _T_261 = io_din[13] & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_262 = _T_258 | _T_261; // @[ifu_compress_ctl.scala 31:22]
  wire  _T_265 = io_din[13] & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_266 = _T_262 | _T_265; // @[ifu_compress_ctl.scala 31:42]
  wire  _T_271 = _T_266 | _T_228; // @[ifu_compress_ctl.scala 31:62]
  wire  out_5 = _T_271 | _T_200; // @[ifu_compress_ctl.scala 31:83]
  wire  _T_288 = _T_2 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_289 = _T_288 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_290 = _T_289 & _T_40; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_291 = _T_290 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_292 = _T_291 & _T_44; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_295 = _T_292 & _T_147; // @[ifu_compress_ctl.scala 33:50]
  wire  _T_303 = _T_194 & _T_147; // @[ifu_compress_ctl.scala 33:87]
  wire  _T_304 = _T_295 | _T_303; // @[ifu_compress_ctl.scala 33:65]
  wire  _T_308 = _T_2 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_311 = _T_308 & _T_147; // @[ifu_compress_ctl.scala 34:23]
  wire  _T_312 = _T_304 | _T_311; // @[ifu_compress_ctl.scala 33:102]
  wire  _T_317 = _T_190 & io_din[14]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_318 = _T_317 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_319 = _T_312 | _T_318; // @[ifu_compress_ctl.scala 34:38]
  wire  _T_323 = _T_2 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_326 = _T_323 & _T_147; // @[ifu_compress_ctl.scala 34:82]
  wire  _T_327 = _T_319 | _T_326; // @[ifu_compress_ctl.scala 34:62]
  wire  _T_331 = _T_2 & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_334 = _T_331 & _T_147; // @[ifu_compress_ctl.scala 35:23]
  wire  _T_335 = _T_327 | _T_334; // @[ifu_compress_ctl.scala 34:97]
  wire  _T_339 = _T_2 & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_342 = _T_339 & _T_147; // @[ifu_compress_ctl.scala 35:58]
  wire  _T_343 = _T_335 | _T_342; // @[ifu_compress_ctl.scala 35:38]
  wire  _T_347 = _T_2 & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_350 = _T_347 & _T_147; // @[ifu_compress_ctl.scala 35:93]
  wire  _T_351 = _T_343 | _T_350; // @[ifu_compress_ctl.scala 35:73]
  wire  _T_357 = _T_2 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_358 = _T_357 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_4 = _T_351 | _T_358; // @[ifu_compress_ctl.scala 35:108]
  wire  _T_380 = _T_56 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_381 = _T_380 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_382 = _T_381 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_383 = _T_382 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_384 = _T_383 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_385 = _T_384 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_386 = _T_385 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_403 = _T_56 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_404 = _T_403 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_405 = _T_404 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_406 = _T_405 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_407 = _T_406 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_408 = _T_407 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_409 = _T_408 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_410 = _T_386 | _T_409; // @[ifu_compress_ctl.scala 40:59]
  wire  _T_427 = _T_56 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_428 = _T_427 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_429 = _T_428 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_430 = _T_429 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_431 = _T_430 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_432 = _T_431 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_433 = _T_432 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_434 = _T_410 | _T_433; // @[ifu_compress_ctl.scala 40:107]
  wire  _T_451 = _T_56 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_452 = _T_451 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_453 = _T_452 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_454 = _T_453 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_455 = _T_454 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_456 = _T_455 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_457 = _T_456 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_458 = _T_434 | _T_457; // @[ifu_compress_ctl.scala 41:50]
  wire  _T_475 = _T_56 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_476 = _T_475 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_477 = _T_476 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_478 = _T_477 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_479 = _T_478 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_480 = _T_479 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_481 = _T_480 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_482 = _T_458 | _T_481; // @[ifu_compress_ctl.scala 41:94]
  wire  _T_487 = ~io_din[12]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_499 = _T_11 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_500 = _T_499 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_501 = _T_500 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_502 = _T_501 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_503 = _T_502 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_504 = _T_503 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_507 = _T_504 & _T_147; // @[ifu_compress_ctl.scala 42:94]
  wire  _T_508 = _T_482 | _T_507; // @[ifu_compress_ctl.scala 42:49]
  wire  _T_514 = _T_190 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_515 = _T_514 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_516 = _T_508 | _T_515; // @[ifu_compress_ctl.scala 42:109]
  wire  _T_522 = _T_514 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_523 = _T_516 | _T_522; // @[ifu_compress_ctl.scala 43:26]
  wire  _T_529 = _T_514 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_530 = _T_523 | _T_529; // @[ifu_compress_ctl.scala 43:48]
  wire  _T_536 = _T_514 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_537 = _T_530 | _T_536; // @[ifu_compress_ctl.scala 43:70]
  wire  _T_543 = _T_514 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_544 = _T_537 | _T_543; // @[ifu_compress_ctl.scala 43:93]
  wire  out_2 = _T_544 | _T_228; // @[ifu_compress_ctl.scala 44:26]
  wire [4:0] rs2d = io_din[6:2]; // @[ifu_compress_ctl.scala 50:20]
  wire [4:0] rdd = io_din[11:7]; // @[ifu_compress_ctl.scala 51:19]
  wire [4:0] rdpd = {2'h1,io_din[9:7]}; // @[Cat.scala 29:58]
  wire [4:0] rs2pd = {2'h1,io_din[4:2]}; // @[Cat.scala 29:58]
  wire  _T_557 = _T_308 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_564 = _T_317 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_565 = _T_564 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_566 = _T_557 | _T_565; // @[ifu_compress_ctl.scala 55:33]
  wire  _T_572 = _T_323 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_573 = _T_566 | _T_572; // @[ifu_compress_ctl.scala 55:58]
  wire  _T_580 = _T_317 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_581 = _T_580 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_582 = _T_573 | _T_581; // @[ifu_compress_ctl.scala 55:79]
  wire  _T_588 = _T_331 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_589 = _T_582 | _T_588; // @[ifu_compress_ctl.scala 55:104]
  wire  _T_596 = _T_317 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_597 = _T_596 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_598 = _T_589 | _T_597; // @[ifu_compress_ctl.scala 56:24]
  wire  _T_604 = _T_339 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_605 = _T_598 | _T_604; // @[ifu_compress_ctl.scala 56:48]
  wire  _T_613 = _T_317 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_614 = _T_613 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_615 = _T_605 | _T_614; // @[ifu_compress_ctl.scala 56:69]
  wire  _T_621 = _T_347 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_622 = _T_615 | _T_621; // @[ifu_compress_ctl.scala 56:94]
  wire  _T_629 = _T_317 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_630 = _T_629 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_631 = _T_622 | _T_630; // @[ifu_compress_ctl.scala 57:22]
  wire  _T_635 = _T_190 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_636 = _T_631 | _T_635; // @[ifu_compress_ctl.scala 57:46]
  wire  _T_642 = _T_190 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_643 = _T_642 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  rdrd = _T_636 | _T_643; // @[ifu_compress_ctl.scala 57:65]
  wire  _T_651 = _T_380 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_659 = _T_403 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_660 = _T_651 | _T_659; // @[ifu_compress_ctl.scala 59:38]
  wire  _T_668 = _T_427 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_669 = _T_660 | _T_668; // @[ifu_compress_ctl.scala 59:63]
  wire  _T_677 = _T_451 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_678 = _T_669 | _T_677; // @[ifu_compress_ctl.scala 59:87]
  wire  _T_686 = _T_475 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_687 = _T_678 | _T_686; // @[ifu_compress_ctl.scala 60:27]
  wire  _T_703 = _T_2 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_704 = _T_703 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_705 = _T_704 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_706 = _T_705 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_707 = _T_706 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_708 = _T_707 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_709 = _T_708 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_710 = _T_687 | _T_709; // @[ifu_compress_ctl.scala 60:51]
  wire  _T_717 = _T_56 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_718 = _T_717 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_719 = _T_710 | _T_718; // @[ifu_compress_ctl.scala 60:89]
  wire  _T_726 = _T_56 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_727 = _T_726 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_728 = _T_719 | _T_727; // @[ifu_compress_ctl.scala 61:27]
  wire  _T_735 = _T_56 & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_736 = _T_735 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_737 = _T_728 | _T_736; // @[ifu_compress_ctl.scala 61:51]
  wire  _T_744 = _T_56 & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_745 = _T_744 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_746 = _T_737 | _T_745; // @[ifu_compress_ctl.scala 61:75]
  wire  _T_753 = _T_56 & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_754 = _T_753 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_755 = _T_746 | _T_754; // @[ifu_compress_ctl.scala 61:99]
  wire  _T_764 = _T_194 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_765 = _T_764 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_766 = _T_755 | _T_765; // @[ifu_compress_ctl.scala 62:27]
  wire  rdrs1 = _T_766 | _T_195; // @[ifu_compress_ctl.scala 62:54]
  wire  _T_777 = io_din[15] & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_778 = _T_777 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_782 = io_din[15] & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_783 = _T_782 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_784 = _T_778 | _T_783; // @[ifu_compress_ctl.scala 64:34]
  wire  _T_788 = io_din[15] & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_789 = _T_788 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_790 = _T_784 | _T_789; // @[ifu_compress_ctl.scala 64:54]
  wire  _T_794 = io_din[15] & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_795 = _T_794 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_796 = _T_790 | _T_795; // @[ifu_compress_ctl.scala 64:74]
  wire  _T_800 = io_din[15] & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_801 = _T_800 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_802 = _T_796 | _T_801; // @[ifu_compress_ctl.scala 64:94]
  wire  _T_807 = _T_200 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  rs2rs2 = _T_802 | _T_807; // @[ifu_compress_ctl.scala 64:114]
  wire  rdprd = _T_12 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_820 = io_din[15] & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_821 = _T_820 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_827 = _T_821 | _T_234; // @[ifu_compress_ctl.scala 68:36]
  wire  _T_830 = ~io_din[1]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_831 = io_din[14] & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_834 = _T_831 & _T_147; // @[ifu_compress_ctl.scala 68:76]
  wire  rdprs1 = _T_827 | _T_834; // @[ifu_compress_ctl.scala 68:57]
  wire  _T_846 = _T_128 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_847 = _T_846 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_851 = io_din[15] & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_854 = _T_851 & _T_147; // @[ifu_compress_ctl.scala 70:66]
  wire  rs2prs2 = _T_847 | _T_854; // @[ifu_compress_ctl.scala 70:47]
  wire  _T_859 = _T_190 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  rs2prd = _T_859 & _T_147; // @[ifu_compress_ctl.scala 72:33]
  wire  _T_866 = _T_2 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  uimm9_2 = _T_866 & _T_147; // @[ifu_compress_ctl.scala 74:34]
  wire  _T_875 = _T_317 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  ulwimm6_2 = _T_875 & _T_147; // @[ifu_compress_ctl.scala 76:39]
  wire  ulwspimm7_2 = _T_317 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_897 = _T_317 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_898 = _T_897 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_899 = _T_898 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_900 = _T_899 & _T_40; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_901 = _T_900 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  rdeq2 = _T_901 & _T_44; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1027 = _T_194 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  rdeq1 = _T_482 | _T_1027; // @[ifu_compress_ctl.scala 84:42]
  wire  _T_1050 = io_din[14] & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1051 = rdeq2 | _T_1050; // @[ifu_compress_ctl.scala 86:53]
  wire  rs1eq2 = _T_1051 | uimm9_2; // @[ifu_compress_ctl.scala 86:71]
  wire  _T_1092 = _T_357 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1093 = _T_1092 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1094 = _T_1093 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  simm5_0 = _T_1094 | _T_643; // @[ifu_compress_ctl.scala 92:45]
  wire  _T_1112 = _T_897 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1121 = _T_897 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1122 = _T_1112 | _T_1121; // @[ifu_compress_ctl.scala 96:44]
  wire  _T_1130 = _T_897 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1131 = _T_1122 | _T_1130; // @[ifu_compress_ctl.scala 96:70]
  wire  _T_1139 = _T_897 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1140 = _T_1131 | _T_1139; // @[ifu_compress_ctl.scala 96:95]
  wire  _T_1148 = _T_897 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  sluimm17_12 = _T_1140 | _T_1148; // @[ifu_compress_ctl.scala 96:121]
  wire  uimm5_0 = _T_79 | _T_195; // @[ifu_compress_ctl.scala 98:45]
  wire [6:0] l1_6 = {out_6,out_5,out_4,_T_228,out_2,1'h1,1'h1}; // @[Cat.scala 29:58]
  wire [4:0] _T_1192 = rdrd ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1193 = rdprd ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1194 = rs2prd ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1195 = rdeq1 ? 5'h1 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1196 = rdeq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1197 = _T_1192 | _T_1193; // @[Mux.scala 27:72]
  wire [4:0] _T_1198 = _T_1197 | _T_1194; // @[Mux.scala 27:72]
  wire [4:0] _T_1199 = _T_1198 | _T_1195; // @[Mux.scala 27:72]
  wire [4:0] l1_11 = _T_1199 | _T_1196; // @[Mux.scala 27:72]
  wire [4:0] _T_1210 = rdrs1 ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1211 = rdprs1 ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1212 = rs1eq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1213 = _T_1210 | _T_1211; // @[Mux.scala 27:72]
  wire [4:0] l1_19 = _T_1213 | _T_1212; // @[Mux.scala 27:72]
  wire [4:0] _T_1219 = {3'h0,1'h0,out_20}; // @[Cat.scala 29:58]
  wire [4:0] _T_1222 = rs2rs2 ? rs2d : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1223 = rs2prs2 ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1224 = _T_1222 | _T_1223; // @[Mux.scala 27:72]
  wire [4:0] l1_24 = _T_1219 | _T_1224; // @[ifu_compress_ctl.scala 114:67]
  wire [14:0] _T_1232 = {out_14,out_13,out_12,l1_11,l1_6}; // @[Cat.scala 29:58]
  wire [31:0] l1 = {1'h0,out_30,2'h0,3'h0,l1_24,l1_19,_T_1232}; // @[Cat.scala 29:58]
  wire [5:0] simm5d = {io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [5:0] simm9d = {io_din[12],io_din[4:3],io_din[5],io_din[2],io_din[6]}; // @[Cat.scala 29:58]
  wire [10:0] sjald_1 = {io_din[12],io_din[8],io_din[10:9],io_din[6],io_din[7],io_din[2],io_din[11],io_din[5:4],io_din[3]}; // @[Cat.scala 29:58]
  wire [19:0] sjald = {io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],sjald_1}; // @[Cat.scala 29:58]
  wire [9:0] _T_1296 = {io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12]}; // @[Cat.scala 29:58]
  wire [19:0] sluimmd = {_T_1296,io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [11:0] _T_1314 = {simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[4:0]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1317 = {2'h0,io_din[10:7],io_din[12:11],io_din[5],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1325 = {simm9d[5],simm9d[5],simm9d[5],simm9d[4:0],4'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1328 = {5'h0,io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1331 = {4'h0,io_din[3:2],io_din[12],io_din[6:4],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1333 = {6'h0,io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [11:0] _T_1339 = {sjald[19],sjald[9:0],sjald[10]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1342 = simm5_0 ? _T_1314 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1343 = uimm9_2 ? _T_1317 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1344 = rdeq2 ? _T_1325 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1345 = ulwimm6_2 ? _T_1328 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1346 = ulwspimm7_2 ? _T_1331 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1347 = uimm5_0 ? _T_1333 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1348 = _T_228 ? _T_1339 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1349 = sluimm17_12 ? sluimmd[19:8] : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1350 = _T_1342 | _T_1343; // @[Mux.scala 27:72]
  wire [11:0] _T_1351 = _T_1350 | _T_1344; // @[Mux.scala 27:72]
  wire [11:0] _T_1352 = _T_1351 | _T_1345; // @[Mux.scala 27:72]
  wire [11:0] _T_1353 = _T_1352 | _T_1346; // @[Mux.scala 27:72]
  wire [11:0] _T_1354 = _T_1353 | _T_1347; // @[Mux.scala 27:72]
  wire [11:0] _T_1355 = _T_1354 | _T_1348; // @[Mux.scala 27:72]
  wire [11:0] _T_1356 = _T_1355 | _T_1349; // @[Mux.scala 27:72]
  wire [11:0] l2_31 = l1[31:20] | _T_1356; // @[ifu_compress_ctl.scala 133:25]
  wire [7:0] _T_1363 = _T_228 ? sjald[19:12] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1364 = sluimm17_12 ? sluimmd[7:0] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1365 = _T_1363 | _T_1364; // @[Mux.scala 27:72]
  wire [7:0] l2_19 = l1[19:12] | _T_1365; // @[ifu_compress_ctl.scala 143:25]
  wire [31:0] l2 = {l2_31,l2_19,l1[11:0]}; // @[Cat.scala 29:58]
  wire [8:0] sbr8d = {io_din[12],io_din[6],io_din[5],io_din[2],io_din[11],io_din[10],io_din[4],io_din[3],1'h0}; // @[Cat.scala 29:58]
  wire [6:0] uswimm6d = {io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [7:0] uswspimm7d = {io_din[8:7],io_din[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [6:0] _T_1400 = {sbr8d[8],sbr8d[8],sbr8d[8],sbr8d[8],sbr8d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1403 = {5'h0,uswimm6d[6:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1406 = {4'h0,uswspimm7d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1407 = _T_234 ? _T_1400 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1408 = _T_854 ? _T_1403 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1409 = _T_807 ? _T_1406 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1410 = _T_1407 | _T_1408; // @[Mux.scala 27:72]
  wire [6:0] _T_1411 = _T_1410 | _T_1409; // @[Mux.scala 27:72]
  wire [6:0] l3_31 = l2[31:25] | _T_1411; // @[ifu_compress_ctl.scala 151:25]
  wire [12:0] l3_24 = l2[24:12]; // @[ifu_compress_ctl.scala 154:17]
  wire [4:0] _T_1417 = {sbr8d[4:1],sbr8d[8]}; // @[Cat.scala 29:58]
  wire [4:0] _T_1422 = _T_234 ? _T_1417 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1423 = _T_854 ? uswimm6d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1424 = _T_807 ? uswspimm7d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1425 = _T_1422 | _T_1423; // @[Mux.scala 27:72]
  wire [4:0] _T_1426 = _T_1425 | _T_1424; // @[Mux.scala 27:72]
  wire [4:0] l3_11 = l2[11:7] | _T_1426; // @[ifu_compress_ctl.scala 156:24]
  wire [31:0] l3 = {l3_31,l3_24,l3_11,l2[6:0]}; // @[Cat.scala 29:58]
  wire  _T_1437 = _T_4 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1438 = _T_1437 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1439 = _T_1438 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1442 = _T_1439 & _T_147; // @[ifu_compress_ctl.scala 162:39]
  wire  _T_1450 = _T_1437 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1451 = _T_1450 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1454 = _T_1451 & _T_147; // @[ifu_compress_ctl.scala 162:79]
  wire  _T_1455 = _T_1442 | _T_1454; // @[ifu_compress_ctl.scala 162:54]
  wire  _T_1464 = _T_642 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1465 = _T_1464 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1466 = _T_1455 | _T_1465; // @[ifu_compress_ctl.scala 162:94]
  wire  _T_1474 = _T_1437 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1475 = _T_1474 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1478 = _T_1475 & _T_147; // @[ifu_compress_ctl.scala 163:55]
  wire  _T_1479 = _T_1466 | _T_1478; // @[ifu_compress_ctl.scala 163:30]
  wire  _T_1487 = _T_1437 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1488 = _T_1487 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1491 = _T_1488 & _T_147; // @[ifu_compress_ctl.scala 163:96]
  wire  _T_1492 = _T_1479 | _T_1491; // @[ifu_compress_ctl.scala 163:70]
  wire  _T_1501 = _T_642 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1502 = _T_1501 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1503 = _T_1492 | _T_1502; // @[ifu_compress_ctl.scala 163:111]
  wire  _T_1510 = io_din[15] & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1511 = _T_1510 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1512 = _T_1511 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1513 = _T_1503 | _T_1512; // @[ifu_compress_ctl.scala 164:29]
  wire  _T_1521 = _T_1437 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1522 = _T_1521 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1525 = _T_1522 & _T_147; // @[ifu_compress_ctl.scala 164:79]
  wire  _T_1526 = _T_1513 | _T_1525; // @[ifu_compress_ctl.scala 164:54]
  wire  _T_1533 = _T_487 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1534 = _T_1533 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1535 = _T_1534 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1536 = _T_1526 | _T_1535; // @[ifu_compress_ctl.scala 164:94]
  wire  _T_1545 = _T_642 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1546 = _T_1545 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1547 = _T_1536 | _T_1546; // @[ifu_compress_ctl.scala 164:118]
  wire  _T_1555 = _T_1437 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1556 = _T_1555 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1559 = _T_1556 & _T_147; // @[ifu_compress_ctl.scala 165:28]
  wire  _T_1560 = _T_1547 | _T_1559; // @[ifu_compress_ctl.scala 164:144]
  wire  _T_1567 = _T_487 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1568 = _T_1567 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1569 = _T_1568 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1570 = _T_1560 | _T_1569; // @[ifu_compress_ctl.scala 165:43]
  wire  _T_1579 = _T_642 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1580 = _T_1579 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1581 = _T_1570 | _T_1580; // @[ifu_compress_ctl.scala 165:67]
  wire  _T_1589 = _T_1437 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1590 = _T_1589 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1593 = _T_1590 & _T_147; // @[ifu_compress_ctl.scala 166:28]
  wire  _T_1594 = _T_1581 | _T_1593; // @[ifu_compress_ctl.scala 165:94]
  wire  _T_1602 = io_din[12] & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1603 = _T_1602 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1604 = _T_1603 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1605 = _T_1604 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1606 = _T_1594 | _T_1605; // @[ifu_compress_ctl.scala 166:43]
  wire  _T_1615 = _T_642 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1616 = _T_1615 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1617 = _T_1606 | _T_1616; // @[ifu_compress_ctl.scala 166:71]
  wire  _T_1625 = _T_1437 & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1626 = _T_1625 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1629 = _T_1626 & _T_147; // @[ifu_compress_ctl.scala 167:28]
  wire  _T_1630 = _T_1617 | _T_1629; // @[ifu_compress_ctl.scala 166:97]
  wire  _T_1636 = io_din[13] & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1637 = _T_1636 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1638 = _T_1637 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1639 = _T_1630 | _T_1638; // @[ifu_compress_ctl.scala 167:43]
  wire  _T_1648 = _T_642 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1649 = _T_1648 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1650 = _T_1639 | _T_1649; // @[ifu_compress_ctl.scala 167:67]
  wire  _T_1658 = _T_1437 & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1659 = _T_1658 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1662 = _T_1659 & _T_147; // @[ifu_compress_ctl.scala 168:28]
  wire  _T_1663 = _T_1650 | _T_1662; // @[ifu_compress_ctl.scala 167:93]
  wire  _T_1669 = io_din[13] & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1670 = _T_1669 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1671 = _T_1670 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1672 = _T_1663 | _T_1671; // @[ifu_compress_ctl.scala 168:43]
  wire  _T_1680 = _T_1437 & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1681 = _T_1680 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1684 = _T_1681 & _T_147; // @[ifu_compress_ctl.scala 168:91]
  wire  _T_1685 = _T_1672 | _T_1684; // @[ifu_compress_ctl.scala 168:66]
  wire  _T_1694 = _T_642 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1695 = _T_1694 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1696 = _T_1685 | _T_1695; // @[ifu_compress_ctl.scala 168:106]
  wire  _T_1702 = io_din[13] & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1703 = _T_1702 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1704 = _T_1703 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1705 = _T_1696 | _T_1704; // @[ifu_compress_ctl.scala 169:29]
  wire  _T_1711 = io_din[13] & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1712 = _T_1711 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1713 = _T_1712 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1714 = _T_1705 | _T_1713; // @[ifu_compress_ctl.scala 169:52]
  wire  _T_1720 = io_din[14] & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1721 = _T_1720 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1722 = _T_1714 | _T_1721; // @[ifu_compress_ctl.scala 169:75]
  wire  _T_1731 = _T_703 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1732 = _T_1731 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1733 = _T_1722 | _T_1732; // @[ifu_compress_ctl.scala 169:98]
  wire  _T_1740 = _T_820 & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1741 = _T_1740 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1744 = _T_1741 & _T_147; // @[ifu_compress_ctl.scala 170:54]
  wire  _T_1745 = _T_1733 | _T_1744; // @[ifu_compress_ctl.scala 170:29]
  wire  _T_1754 = _T_642 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1755 = _T_1754 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1758 = _T_1755 & _T_147; // @[ifu_compress_ctl.scala 170:96]
  wire  _T_1759 = _T_1745 | _T_1758; // @[ifu_compress_ctl.scala 170:69]
  wire  _T_1768 = _T_642 & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1769 = _T_1768 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1770 = _T_1759 | _T_1769; // @[ifu_compress_ctl.scala 170:111]
  wire  _T_1777 = _T_1720 & _T_147; // @[ifu_compress_ctl.scala 171:50]
  wire  legal = _T_1770 | _T_1777; // @[ifu_compress_ctl.scala 171:30]
  wire [9:0] _T_1787 = {legal,legal,legal,legal,legal,legal,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  wire [18:0] _T_1796 = {_T_1787,legal,legal,legal,legal,legal,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  wire [27:0] _T_1805 = {_T_1796,legal,legal,legal,legal,legal,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  wire [31:0] _T_1809 = {_T_1805,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  assign io_dout = l3 & _T_1809; // @[ifu_compress_ctl.scala 173:10]
endmodule
module ifu_aln_ctl(
  input         clk,
  input         reset,
  input         io_active_clk,
  input         io_ifu_async_error_start,
  input  [1:0]  io_iccm_rd_ecc_double_err,
  input  [1:0]  io_ic_access_fault_f,
  input  [1:0]  io_ic_access_fault_type_f,
  input         io_dec_i0_decode_d,
  output [15:0] io_dec_aln_aln_dec_ifu_i0_cinst,
  output        io_dec_aln_aln_ib_ifu_i0_icaf,
  output [1:0]  io_dec_aln_aln_ib_ifu_i0_icaf_type,
  output        io_dec_aln_aln_ib_ifu_i0_icaf_second,
  output        io_dec_aln_aln_ib_ifu_i0_dbecc,
  output [7:0]  io_dec_aln_aln_ib_ifu_i0_bp_index,
  output [7:0]  io_dec_aln_aln_ib_ifu_i0_bp_fghr,
  output [4:0]  io_dec_aln_aln_ib_ifu_i0_bp_btag,
  output        io_dec_aln_aln_ib_ifu_i0_valid,
  output [31:0] io_dec_aln_aln_ib_ifu_i0_instr,
  output [30:0] io_dec_aln_aln_ib_ifu_i0_pc,
  output        io_dec_aln_aln_ib_ifu_i0_pc4,
  output        io_dec_aln_aln_ib_i0_brp_valid,
  output [11:0] io_dec_aln_aln_ib_i0_brp_bits_toffset,
  output [1:0]  io_dec_aln_aln_ib_i0_brp_bits_hist,
  output        io_dec_aln_aln_ib_i0_brp_bits_br_error,
  output        io_dec_aln_aln_ib_i0_brp_bits_br_start_error,
  output        io_dec_aln_aln_ib_i0_brp_bits_bank,
  output [30:0] io_dec_aln_aln_ib_i0_brp_bits_prett,
  output        io_dec_aln_aln_ib_i0_brp_bits_way,
  output        io_dec_aln_aln_ib_i0_brp_bits_ret,
  output        io_dec_aln_ifu_pmu_instr_aligned,
  input  [7:0]  io_ifu_bp_fghr_f,
  input  [30:0] io_ifu_bp_btb_target_f,
  input  [11:0] io_ifu_bp_poffset_f,
  input  [1:0]  io_ifu_bp_hist0_f,
  input  [1:0]  io_ifu_bp_hist1_f,
  input  [1:0]  io_ifu_bp_pc4_f,
  input  [1:0]  io_ifu_bp_way_f,
  input  [1:0]  io_ifu_bp_valid_f,
  input  [1:0]  io_ifu_bp_ret_f,
  input         io_exu_flush_final,
  input  [31:0] io_ifu_fetch_data_f,
  input  [1:0]  io_ifu_fetch_val,
  input  [30:0] io_ifu_fetch_pc,
  output        io_ifu_fb_consume1,
  output        io_ifu_fb_consume2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 409:23]
  wire [15:0] decompressed_io_din; // @[ifu_aln_ctl.scala 444:28]
  wire [31:0] decompressed_io_dout; // @[ifu_aln_ctl.scala 444:28]
  reg  error_stall; // @[Reg.scala 27:20]
  wire  _T = error_stall | io_ifu_async_error_start; // @[ifu_aln_ctl.scala 119:37]
  wire  _T_1 = ~io_exu_flush_final; // @[ifu_aln_ctl.scala 119:67]
  wire  error_stall_in = _T & _T_1; // @[ifu_aln_ctl.scala 119:65]
  reg [1:0] wrptr; // @[ifu_aln_ctl.scala 120:48]
  reg [1:0] rdptr; // @[ifu_aln_ctl.scala 121:48]
  reg  q2off; // @[ifu_aln_ctl.scala 122:48]
  reg  q1off; // @[ifu_aln_ctl.scala 123:48]
  reg  q0off; // @[ifu_aln_ctl.scala 124:48]
  wire  _T_3 = error_stall_in ^ error_stall; // @[lib.scala 453:21]
  wire  _T_4 = |_T_3; // @[lib.scala 453:29]
  wire  _T_821 = ~error_stall; // @[ifu_aln_ctl.scala 504:39]
  wire  i0_shift = io_dec_i0_decode_d & _T_821; // @[ifu_aln_ctl.scala 504:37]
  reg [1:0] f0val; // @[Reg.scala 27:20]
  wire  _T_191 = rdptr == 2'h0; // @[ifu_aln_ctl.scala 192:31]
  wire  _T_194 = _T_191 & q0off; // @[Mux.scala 27:72]
  wire  _T_192 = rdptr == 2'h1; // @[ifu_aln_ctl.scala 193:11]
  wire  _T_195 = _T_192 & q1off; // @[Mux.scala 27:72]
  wire  _T_197 = _T_194 | _T_195; // @[Mux.scala 27:72]
  wire  _T_193 = rdptr == 2'h2; // @[ifu_aln_ctl.scala 194:11]
  wire  _T_196 = _T_193 & q2off; // @[Mux.scala 27:72]
  wire  q0ptr = _T_197 | _T_196; // @[Mux.scala 27:72]
  wire  _T_207 = ~q0ptr; // @[ifu_aln_ctl.scala 198:26]
  wire [1:0] q0sel = {q0ptr,_T_207}; // @[Cat.scala 29:58]
  wire [2:0] qren = {_T_193,_T_192,_T_191}; // @[Cat.scala 29:58]
  reg [31:0] q1; // @[Reg.scala 27:20]
  reg [31:0] q0; // @[Reg.scala 27:20]
  wire [63:0] _T_479 = {q1,q0}; // @[Cat.scala 29:58]
  wire [63:0] _T_486 = qren[0] ? _T_479 : 64'h0; // @[Mux.scala 27:72]
  reg [31:0] q2; // @[Reg.scala 27:20]
  wire [63:0] _T_482 = {q2,q1}; // @[Cat.scala 29:58]
  wire [63:0] _T_487 = qren[1] ? _T_482 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_489 = _T_486 | _T_487; // @[Mux.scala 27:72]
  wire [63:0] _T_485 = {q0,q2}; // @[Cat.scala 29:58]
  wire [63:0] _T_488 = qren[2] ? _T_485 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] qeff = _T_489 | _T_488; // @[Mux.scala 27:72]
  wire [31:0] q0eff = qeff[31:0]; // @[ifu_aln_ctl.scala 370:42]
  wire [31:0] _T_496 = q0sel[0] ? q0eff : 32'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_497 = q0sel[1] ? q0eff[31:16] : 16'h0; // @[Mux.scala 27:72]
  wire [31:0] _GEN_16 = {{16'd0}, _T_497}; // @[Mux.scala 27:72]
  wire [31:0] q0final = _T_496 | _GEN_16; // @[Mux.scala 27:72]
  wire [31:0] _T_541 = f0val[1] ? q0final : 32'h0; // @[Mux.scala 27:72]
  wire  _T_534 = ~f0val[1]; // @[ifu_aln_ctl.scala 384:58]
  wire  _T_536 = _T_534 & f0val[0]; // @[ifu_aln_ctl.scala 384:68]
  wire  _T_202 = _T_191 & q1off; // @[Mux.scala 27:72]
  wire  _T_203 = _T_192 & q2off; // @[Mux.scala 27:72]
  wire  _T_205 = _T_202 | _T_203; // @[Mux.scala 27:72]
  wire  _T_204 = _T_193 & q0off; // @[Mux.scala 27:72]
  wire  q1ptr = _T_205 | _T_204; // @[Mux.scala 27:72]
  wire  _T_208 = ~q1ptr; // @[ifu_aln_ctl.scala 200:26]
  wire [1:0] q1sel = {q1ptr,_T_208}; // @[Cat.scala 29:58]
  wire [31:0] q1eff = qeff[63:32]; // @[ifu_aln_ctl.scala 370:29]
  wire [15:0] _T_506 = q1sel[0] ? q1eff[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_507 = q1sel[1] ? q1eff[31:16] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] q1final = _T_506 | _T_507; // @[Mux.scala 27:72]
  wire [31:0] _T_540 = {q1final,q0final[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_542 = _T_536 ? _T_540 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] aligndata = _T_541 | _T_542; // @[Mux.scala 27:72]
  wire  first4B = aligndata[1:0] == 2'h3; // @[ifu_aln_ctl.scala 426:29]
  wire  first2B = ~first4B; // @[ifu_aln_ctl.scala 428:17]
  wire  shift_2B = i0_shift & first2B; // @[ifu_aln_ctl.scala 508:24]
  wire [1:0] _T_443 = {1'h0,f0val[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_448 = shift_2B ? _T_443 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_444 = ~shift_2B; // @[ifu_aln_ctl.scala 360:6]
  wire  shift_4B = i0_shift & first4B; // @[ifu_aln_ctl.scala 509:24]
  wire  _T_445 = ~shift_4B; // @[ifu_aln_ctl.scala 360:18]
  wire  _T_446 = _T_444 & _T_445; // @[ifu_aln_ctl.scala 360:16]
  wire [1:0] _T_449 = _T_446 ? f0val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] sf0val = _T_448 | _T_449; // @[Mux.scala 27:72]
  wire  sf0_valid = sf0val[0]; // @[ifu_aln_ctl.scala 326:22]
  wire  _T_389 = ~sf0_valid; // @[ifu_aln_ctl.scala 347:26]
  wire  _T_838 = f0val[0] & _T_534; // @[ifu_aln_ctl.scala 512:28]
  wire  f1_shift_2B = _T_838 & shift_4B; // @[ifu_aln_ctl.scala 512:40]
  reg [1:0] f1val; // @[Reg.scala 27:20]
  wire  _T_417 = f1_shift_2B & f1val[1]; // @[Mux.scala 27:72]
  wire  _T_416 = ~f1_shift_2B; // @[ifu_aln_ctl.scala 353:53]
  wire [1:0] _T_418 = _T_416 ? f1val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_17 = {{1'd0}, _T_417}; // @[Mux.scala 27:72]
  wire [1:0] sf1val = _GEN_17 | _T_418; // @[Mux.scala 27:72]
  wire  sf1_valid = sf1val[0]; // @[ifu_aln_ctl.scala 325:22]
  wire  _T_390 = _T_389 & sf1_valid; // @[ifu_aln_ctl.scala 347:37]
  reg [1:0] f2val; // @[Reg.scala 27:20]
  wire  f2_valid = f2val[0]; // @[ifu_aln_ctl.scala 324:20]
  wire  _T_391 = _T_390 & f2_valid; // @[ifu_aln_ctl.scala 347:50]
  wire  ifvalid = io_ifu_fetch_val[0]; // @[ifu_aln_ctl.scala 335:30]
  wire  _T_392 = _T_391 & ifvalid; // @[ifu_aln_ctl.scala 347:62]
  wire  _T_393 = sf0_valid & sf1_valid; // @[ifu_aln_ctl.scala 348:17]
  wire  _T_394 = ~f2_valid; // @[ifu_aln_ctl.scala 348:32]
  wire  _T_395 = _T_393 & _T_394; // @[ifu_aln_ctl.scala 348:30]
  wire  _T_396 = _T_395 & ifvalid; // @[ifu_aln_ctl.scala 348:42]
  wire  fetch_to_f2 = _T_392 | _T_396; // @[ifu_aln_ctl.scala 347:74]
  wire  _T_399 = fetch_to_f2 & _T_1; // @[ifu_aln_ctl.scala 350:38]
  wire [1:0] _T_409 = _T_399 ? io_ifu_fetch_val : 2'h0; // @[Mux.scala 27:72]
  wire  _T_401 = ~fetch_to_f2; // @[ifu_aln_ctl.scala 351:6]
  wire  _T_402 = ~_T_391; // @[ifu_aln_ctl.scala 351:21]
  wire  _T_403 = _T_401 & _T_402; // @[ifu_aln_ctl.scala 351:19]
  wire  _T_360 = ~sf1_valid; // @[ifu_aln_ctl.scala 339:31]
  wire  _T_361 = _T_389 & _T_360; // @[ifu_aln_ctl.scala 339:29]
  wire  shift_f2_f0 = _T_361 & f2_valid; // @[ifu_aln_ctl.scala 339:42]
  wire  _T_404 = ~shift_f2_f0; // @[ifu_aln_ctl.scala 351:36]
  wire  _T_405 = _T_403 & _T_404; // @[ifu_aln_ctl.scala 351:34]
  wire  _T_407 = _T_405 & _T_1; // @[ifu_aln_ctl.scala 351:49]
  wire [1:0] _T_410 = _T_407 ? f2val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] f2val_in = _T_409 | _T_410; // @[Mux.scala 27:72]
  wire [1:0] _T_6 = f2val_in ^ f2val; // @[lib.scala 453:21]
  wire  _T_7 = |_T_6; // @[lib.scala 453:29]
  wire  _T_376 = shift_f2_f0 & ifvalid; // @[ifu_aln_ctl.scala 343:62]
  wire  _T_380 = _T_390 & _T_394; // @[ifu_aln_ctl.scala 344:30]
  wire  _T_381 = _T_380 & ifvalid; // @[ifu_aln_ctl.scala 344:42]
  wire  _T_382 = _T_376 | _T_381; // @[ifu_aln_ctl.scala 343:74]
  wire  _T_384 = sf0_valid & _T_360; // @[ifu_aln_ctl.scala 345:17]
  wire  _T_386 = _T_384 & _T_394; // @[ifu_aln_ctl.scala 345:30]
  wire  _T_387 = _T_386 & ifvalid; // @[ifu_aln_ctl.scala 345:42]
  wire  fetch_to_f1 = _T_382 | _T_387; // @[ifu_aln_ctl.scala 344:54]
  wire  _T_422 = fetch_to_f1 & _T_1; // @[ifu_aln_ctl.scala 355:39]
  wire [1:0] _T_435 = _T_422 ? io_ifu_fetch_val : 2'h0; // @[Mux.scala 27:72]
  wire  _T_425 = _T_391 & _T_1; // @[ifu_aln_ctl.scala 356:34]
  wire [1:0] _T_436 = _T_425 ? f2val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_438 = _T_435 | _T_436; // @[Mux.scala 27:72]
  wire  _T_427 = ~fetch_to_f1; // @[ifu_aln_ctl.scala 357:6]
  wire  _T_429 = _T_427 & _T_402; // @[ifu_aln_ctl.scala 357:19]
  wire  _T_430 = ~_T_390; // @[ifu_aln_ctl.scala 357:36]
  wire  _T_431 = _T_429 & _T_430; // @[ifu_aln_ctl.scala 357:34]
  wire  _T_433 = _T_431 & _T_1; // @[ifu_aln_ctl.scala 357:49]
  wire [1:0] _T_437 = _T_433 ? sf1val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] f1val_in = _T_438 | _T_437; // @[Mux.scala 27:72]
  wire [1:0] _T_9 = f1val_in ^ f1val; // @[lib.scala 453:21]
  wire  _T_10 = |_T_9; // @[lib.scala 453:29]
  wire  _T_370 = _T_361 & _T_394; // @[ifu_aln_ctl.scala 342:50]
  wire  fetch_to_f0 = _T_370 & ifvalid; // @[ifu_aln_ctl.scala 342:62]
  wire  _T_453 = fetch_to_f0 & _T_1; // @[ifu_aln_ctl.scala 362:38]
  wire [1:0] _T_469 = _T_453 ? io_ifu_fetch_val : 2'h0; // @[Mux.scala 27:72]
  wire  _T_456 = shift_f2_f0 & _T_1; // @[ifu_aln_ctl.scala 363:34]
  wire [1:0] _T_470 = _T_456 ? f2val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_473 = _T_469 | _T_470; // @[Mux.scala 27:72]
  wire  _T_459 = _T_390 & _T_1; // @[ifu_aln_ctl.scala 364:49]
  wire [1:0] _T_471 = _T_459 ? sf1val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_474 = _T_473 | _T_471; // @[Mux.scala 27:72]
  wire  _T_461 = ~fetch_to_f0; // @[ifu_aln_ctl.scala 365:6]
  wire  _T_463 = _T_461 & _T_404; // @[ifu_aln_ctl.scala 365:19]
  wire  _T_465 = _T_463 & _T_430; // @[ifu_aln_ctl.scala 365:34]
  wire  _T_467 = _T_465 & _T_1; // @[ifu_aln_ctl.scala 365:49]
  wire [1:0] _T_472 = _T_467 ? sf0val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] f0val_in = _T_474 | _T_472; // @[Mux.scala 27:72]
  wire [1:0] _T_12 = f0val_in ^ f0val; // @[lib.scala 453:21]
  wire  _T_13 = |_T_12; // @[lib.scala 453:29]
  wire  _T_40 = wrptr == 2'h2; // @[ifu_aln_ctl.scala 162:22]
  wire  _T_41 = _T_40 & ifvalid; // @[ifu_aln_ctl.scala 162:31]
  wire  _T_42 = wrptr == 2'h1; // @[ifu_aln_ctl.scala 162:49]
  wire  _T_43 = _T_42 & ifvalid; // @[ifu_aln_ctl.scala 162:58]
  wire  _T_44 = wrptr == 2'h0; // @[ifu_aln_ctl.scala 162:76]
  wire  _T_45 = _T_44 & ifvalid; // @[ifu_aln_ctl.scala 162:85]
  wire [2:0] qwen = {_T_41,_T_43,_T_45}; // @[Cat.scala 29:58]
  reg [15:0] brdata2; // @[Reg.scala 27:20]
  wire [7:0] _T_283 = {io_iccm_rd_ecc_double_err[0],io_ic_access_fault_f[0],io_ifu_bp_hist1_f[0],io_ifu_bp_hist0_f[0],io_ifu_bp_pc4_f[0],io_ifu_bp_way_f[0],io_ifu_bp_valid_f[0],io_ifu_bp_ret_f[0]}; // @[Cat.scala 29:58]
  wire [15:0] brdata_in = {io_iccm_rd_ecc_double_err[1],io_ic_access_fault_f[1],io_ifu_bp_hist1_f[1],io_ifu_bp_hist0_f[1],io_ifu_bp_pc4_f[1],io_ifu_bp_way_f[1],io_ifu_bp_valid_f[1],io_ifu_bp_ret_f[1],_T_283}; // @[Cat.scala 29:58]
  reg [15:0] brdata1; // @[Reg.scala 27:20]
  reg [15:0] brdata0; // @[Reg.scala 27:20]
  reg [52:0] misc2; // @[Reg.scala 27:20]
  wire [52:0] misc_data_in = {io_ic_access_fault_type_f,io_ifu_bp_btb_target_f,io_ifu_bp_poffset_f,io_ifu_bp_fghr_f}; // @[Cat.scala 29:58]
  reg [52:0] misc1; // @[Reg.scala 27:20]
  reg [52:0] misc0; // @[Reg.scala 27:20]
  reg [30:0] q2pc; // @[Reg.scala 27:20]
  reg [30:0] q1pc; // @[Reg.scala 27:20]
  reg [30:0] q0pc; // @[Reg.scala 27:20]
  wire  _T_49 = qren[0] & io_ifu_fb_consume1; // @[ifu_aln_ctl.scala 164:34]
  wire  _T_51 = _T_49 & _T_1; // @[ifu_aln_ctl.scala 164:55]
  wire  _T_54 = qren[1] & io_ifu_fb_consume1; // @[ifu_aln_ctl.scala 165:14]
  wire  _T_56 = _T_54 & _T_1; // @[ifu_aln_ctl.scala 165:35]
  wire  _T_64 = qren[0] & io_ifu_fb_consume2; // @[ifu_aln_ctl.scala 167:14]
  wire  _T_66 = _T_64 & _T_1; // @[ifu_aln_ctl.scala 167:35]
  wire  _T_74 = qren[2] & io_ifu_fb_consume2; // @[ifu_aln_ctl.scala 169:14]
  wire  _T_76 = _T_74 & _T_1; // @[ifu_aln_ctl.scala 169:35]
  wire  _T_78 = ~io_ifu_fb_consume1; // @[ifu_aln_ctl.scala 170:6]
  wire  _T_79 = ~io_ifu_fb_consume2; // @[ifu_aln_ctl.scala 170:28]
  wire  _T_80 = _T_78 & _T_79; // @[ifu_aln_ctl.scala 170:26]
  wire  _T_82 = _T_80 & _T_1; // @[ifu_aln_ctl.scala 170:48]
  wire [1:0] _T_85 = _T_56 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_87 = _T_66 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_90 = _T_82 ? rdptr : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_18 = {{1'd0}, _T_51}; // @[Mux.scala 27:72]
  wire [1:0] _T_91 = _GEN_18 | _T_85; // @[Mux.scala 27:72]
  wire [1:0] _T_93 = _T_91 | _T_87; // @[Mux.scala 27:72]
  wire [1:0] _GEN_19 = {{1'd0}, _T_76}; // @[Mux.scala 27:72]
  wire [1:0] _T_95 = _T_93 | _GEN_19; // @[Mux.scala 27:72]
  wire  _T_100 = qwen[0] & _T_1; // @[ifu_aln_ctl.scala 173:34]
  wire  _T_104 = qwen[1] & _T_1; // @[ifu_aln_ctl.scala 174:14]
  wire  _T_110 = ~ifvalid; // @[ifu_aln_ctl.scala 176:6]
  wire  _T_112 = _T_110 & _T_1; // @[ifu_aln_ctl.scala 176:15]
  wire [1:0] _T_115 = _T_104 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_117 = _T_112 ? wrptr : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_20 = {{1'd0}, _T_100}; // @[Mux.scala 27:72]
  wire [1:0] _T_118 = _GEN_20 | _T_115; // @[Mux.scala 27:72]
  wire  _T_123 = ~qwen[2]; // @[ifu_aln_ctl.scala 178:26]
  wire  _T_125 = _T_123 & _T_193; // @[ifu_aln_ctl.scala 178:35]
  wire  _T_831 = shift_2B & f0val[0]; // @[Mux.scala 27:72]
  wire  _T_832 = shift_4B & _T_838; // @[Mux.scala 27:72]
  wire  f0_shift_2B = _T_831 | _T_832; // @[Mux.scala 27:72]
  wire  _T_127 = q2off | f0_shift_2B; // @[ifu_aln_ctl.scala 178:76]
  wire  _T_131 = _T_123 & _T_192; // @[ifu_aln_ctl.scala 179:15]
  wire  _T_133 = q2off | f1_shift_2B; // @[ifu_aln_ctl.scala 179:56]
  wire  _T_137 = _T_123 & _T_191; // @[ifu_aln_ctl.scala 180:15]
  wire  _T_139 = _T_125 & _T_127; // @[Mux.scala 27:72]
  wire  _T_140 = _T_131 & _T_133; // @[Mux.scala 27:72]
  wire  _T_141 = _T_137 & q2off; // @[Mux.scala 27:72]
  wire  _T_142 = _T_139 | _T_140; // @[Mux.scala 27:72]
  wire  _T_146 = ~qwen[1]; // @[ifu_aln_ctl.scala 182:26]
  wire  _T_148 = _T_146 & _T_192; // @[ifu_aln_ctl.scala 182:35]
  wire  _T_150 = q1off | f0_shift_2B; // @[ifu_aln_ctl.scala 182:76]
  wire  _T_154 = _T_146 & _T_191; // @[ifu_aln_ctl.scala 183:15]
  wire  _T_156 = q1off | f1_shift_2B; // @[ifu_aln_ctl.scala 183:56]
  wire  _T_160 = _T_146 & _T_193; // @[ifu_aln_ctl.scala 184:15]
  wire  _T_162 = _T_148 & _T_150; // @[Mux.scala 27:72]
  wire  _T_163 = _T_154 & _T_156; // @[Mux.scala 27:72]
  wire  _T_164 = _T_160 & q1off; // @[Mux.scala 27:72]
  wire  _T_165 = _T_162 | _T_163; // @[Mux.scala 27:72]
  wire  _T_169 = ~qwen[0]; // @[ifu_aln_ctl.scala 186:26]
  wire  _T_171 = _T_169 & _T_191; // @[ifu_aln_ctl.scala 186:35]
  wire  _T_173 = q0off | f0_shift_2B; // @[ifu_aln_ctl.scala 186:76]
  wire  _T_177 = _T_169 & _T_193; // @[ifu_aln_ctl.scala 187:15]
  wire  _T_179 = q0off | f1_shift_2B; // @[ifu_aln_ctl.scala 187:56]
  wire  _T_183 = _T_169 & _T_192; // @[ifu_aln_ctl.scala 188:15]
  wire  _T_185 = _T_171 & _T_173; // @[Mux.scala 27:72]
  wire  _T_186 = _T_177 & _T_179; // @[Mux.scala 27:72]
  wire  _T_187 = _T_183 & q0off; // @[Mux.scala 27:72]
  wire  _T_188 = _T_185 | _T_186; // @[Mux.scala 27:72]
  wire [105:0] _T_214 = {misc1,misc0}; // @[Cat.scala 29:58]
  wire [105:0] _T_217 = {misc2,misc1}; // @[Cat.scala 29:58]
  wire [105:0] _T_220 = {misc0,misc2}; // @[Cat.scala 29:58]
  wire [105:0] _T_221 = qren[0] ? _T_214 : 106'h0; // @[Mux.scala 27:72]
  wire [105:0] _T_222 = qren[1] ? _T_217 : 106'h0; // @[Mux.scala 27:72]
  wire [105:0] _T_223 = qren[2] ? _T_220 : 106'h0; // @[Mux.scala 27:72]
  wire [105:0] _T_224 = _T_221 | _T_222; // @[Mux.scala 27:72]
  wire [105:0] misceff = _T_224 | _T_223; // @[Mux.scala 27:72]
  wire [52:0] misc1eff = misceff[105:53]; // @[ifu_aln_ctl.scala 214:25]
  wire [52:0] misc0eff = misceff[52:0]; // @[ifu_aln_ctl.scala 215:25]
  wire [1:0] f1ictype = misc1eff[52:51]; // @[ifu_aln_ctl.scala 218:43]
  wire [30:0] f1prett = misc1eff[50:20]; // @[ifu_aln_ctl.scala 219:43]
  wire [11:0] f1poffset = misc1eff[19:8]; // @[ifu_aln_ctl.scala 220:43]
  wire [7:0] f1fghr = misc1eff[7:0]; // @[ifu_aln_ctl.scala 221:43]
  wire [1:0] f0ictype = misc0eff[52:51]; // @[ifu_aln_ctl.scala 223:43]
  wire [30:0] f0prett = misc0eff[50:20]; // @[ifu_aln_ctl.scala 224:43]
  wire [11:0] f0poffset = misc0eff[19:8]; // @[ifu_aln_ctl.scala 225:43]
  wire [7:0] f0fghr = misc0eff[7:0]; // @[ifu_aln_ctl.scala 226:43]
  wire [31:0] _T_228 = {brdata1,brdata0}; // @[Cat.scala 29:58]
  wire [31:0] _T_231 = {brdata2,brdata1}; // @[Cat.scala 29:58]
  wire [31:0] _T_234 = {brdata0,brdata2}; // @[Cat.scala 29:58]
  wire [31:0] _T_235 = qren[0] ? _T_228 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_236 = qren[1] ? _T_231 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_237 = qren[2] ? _T_234 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_238 = _T_235 | _T_236; // @[Mux.scala 27:72]
  wire [31:0] brdataeff = _T_238 | _T_237; // @[Mux.scala 27:72]
  wire [15:0] brdata1eff = brdataeff[31:16]; // @[ifu_aln_ctl.scala 254:26]
  wire [15:0] brdata0eff = brdataeff[15:0]; // @[ifu_aln_ctl.scala 255:26]
  wire [15:0] _T_249 = q0sel[0] ? brdata0eff : 16'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_250 = q0sel[1] ? brdata0eff[15:8] : 8'h0; // @[Mux.scala 27:72]
  wire [15:0] _GEN_21 = {{8'd0}, _T_250}; // @[Mux.scala 27:72]
  wire [15:0] brdata0final = _T_249 | _GEN_21; // @[Mux.scala 27:72]
  wire [15:0] _T_258 = q1sel[0] ? brdata1eff : 16'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_259 = q1sel[1] ? brdata1eff[15:8] : 8'h0; // @[Mux.scala 27:72]
  wire [15:0] _GEN_22 = {{8'd0}, _T_259}; // @[Mux.scala 27:72]
  wire [15:0] brdata1final = _T_258 | _GEN_22; // @[Mux.scala 27:72]
  wire [1:0] f0ret = {brdata0final[8],brdata0final[0]}; // @[Cat.scala 29:58]
  wire [1:0] f0brend = {brdata0final[9],brdata0final[1]}; // @[Cat.scala 29:58]
  wire [1:0] f0way = {brdata0final[10],brdata0final[2]}; // @[Cat.scala 29:58]
  wire [1:0] f0pc4 = {brdata0final[11],brdata0final[3]}; // @[Cat.scala 29:58]
  wire [1:0] f0hist0 = {brdata0final[12],brdata0final[4]}; // @[Cat.scala 29:58]
  wire [1:0] f0hist1 = {brdata0final[13],brdata0final[5]}; // @[Cat.scala 29:58]
  wire [1:0] f0icaf = {brdata0final[14],brdata0final[6]}; // @[Cat.scala 29:58]
  wire [1:0] f0dbecc = {brdata0final[15],brdata0final[7]}; // @[Cat.scala 29:58]
  wire [1:0] f1ret = {brdata1final[8],brdata1final[0]}; // @[Cat.scala 29:58]
  wire [1:0] f1brend = {brdata1final[9],brdata1final[1]}; // @[Cat.scala 29:58]
  wire [1:0] f1way = {brdata1final[10],brdata1final[2]}; // @[Cat.scala 29:58]
  wire [1:0] f1pc4 = {brdata1final[11],brdata1final[3]}; // @[Cat.scala 29:58]
  wire [1:0] f1hist0 = {brdata1final[12],brdata1final[4]}; // @[Cat.scala 29:58]
  wire [1:0] f1hist1 = {brdata1final[13],brdata1final[5]}; // @[Cat.scala 29:58]
  wire [1:0] f1icaf = {brdata1final[14],brdata1final[6]}; // @[Cat.scala 29:58]
  wire [1:0] f1dbecc = {brdata1final[15],brdata1final[7]}; // @[Cat.scala 29:58]
  wire  consume_fb0 = _T_389 & f0val[0]; // @[ifu_aln_ctl.scala 328:32]
  wire  consume_fb1 = _T_360 & f1val[0]; // @[ifu_aln_ctl.scala 329:32]
  wire  _T_349 = ~consume_fb1; // @[ifu_aln_ctl.scala 332:39]
  wire  _T_350 = consume_fb0 & _T_349; // @[ifu_aln_ctl.scala 332:37]
  wire  _T_353 = consume_fb0 & consume_fb1; // @[ifu_aln_ctl.scala 333:37]
  wire [61:0] _T_512 = {q1pc,q0pc}; // @[Cat.scala 29:58]
  wire [61:0] _T_515 = {q2pc,q1pc}; // @[Cat.scala 29:58]
  wire [61:0] _T_518 = {q0pc,q2pc}; // @[Cat.scala 29:58]
  wire [61:0] _T_519 = qren[0] ? _T_512 : 62'h0; // @[Mux.scala 27:72]
  wire [61:0] _T_520 = qren[1] ? _T_515 : 62'h0; // @[Mux.scala 27:72]
  wire [61:0] _T_521 = qren[2] ? _T_518 : 62'h0; // @[Mux.scala 27:72]
  wire [61:0] _T_522 = _T_519 | _T_520; // @[Mux.scala 27:72]
  wire [61:0] qpceff = _T_522 | _T_521; // @[Mux.scala 27:72]
  wire [30:0] q1pceff = qpceff[61:31]; // @[ifu_aln_ctl.scala 380:23]
  wire [30:0] q0pceff = qpceff[30:0]; // @[ifu_aln_ctl.scala 381:23]
  wire [30:0] _T_527 = q0pceff + 31'h1; // @[ifu_aln_ctl.scala 382:70]
  wire [30:0] _T_528 = q0sel[0] ? q0pceff : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_529 = q0sel[1] ? _T_527 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] firstpc = _T_528 | _T_529; // @[Mux.scala 27:72]
  wire [1:0] _T_551 = {f1val[0],1'h1}; // @[Cat.scala 29:58]
  wire [1:0] _T_552 = f0val[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_553 = _T_536 ? _T_551 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignval = _T_552 | _T_553; // @[Mux.scala 27:72]
  wire [1:0] _T_565 = {f1icaf[0],f0icaf[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_566 = f0val[1] ? f0icaf : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_567 = _T_536 ? _T_565 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignicaf = _T_566 | _T_567; // @[Mux.scala 27:72]
  wire [1:0] _T_578 = {f1dbecc[0],f0dbecc[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_579 = f0val[1] ? f0dbecc : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_580 = _T_536 ? _T_578 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] aligndbecc = _T_579 | _T_580; // @[Mux.scala 27:72]
  wire [1:0] _T_591 = {f1brend[0],f0brend[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_592 = f0val[1] ? f0brend : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_593 = _T_536 ? _T_591 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignbrend = _T_592 | _T_593; // @[Mux.scala 27:72]
  wire [1:0] _T_604 = {f1pc4[0],f0pc4[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_605 = f0val[1] ? f0pc4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_606 = _T_536 ? _T_604 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignpc4 = _T_605 | _T_606; // @[Mux.scala 27:72]
  wire [1:0] _T_617 = {f1ret[0],f0ret[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_618 = f0val[1] ? f0ret : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_619 = _T_536 ? _T_617 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignret = _T_618 | _T_619; // @[Mux.scala 27:72]
  wire [1:0] _T_630 = {f1way[0],f0way[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_631 = f0val[1] ? f0way : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_632 = _T_536 ? _T_630 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignway = _T_631 | _T_632; // @[Mux.scala 27:72]
  wire [1:0] _T_643 = {f1hist1[0],f0hist1[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_644 = f0val[1] ? f0hist1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_645 = _T_536 ? _T_643 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignhist1 = _T_644 | _T_645; // @[Mux.scala 27:72]
  wire [1:0] _T_656 = {f1hist0[0],f0hist0[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_657 = f0val[1] ? f0hist0 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_658 = _T_536 ? _T_656 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignhist0 = _T_657 | _T_658; // @[Mux.scala 27:72]
  wire [30:0] _T_669 = f0val[1] ? _T_527 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_670 = _T_536 ? q1pceff : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] secondpc = _T_669 | _T_670; // @[Mux.scala 27:72]
  wire  _T_682 = first4B & alignval[1]; // @[Mux.scala 27:72]
  wire  _T_683 = first2B & alignval[0]; // @[Mux.scala 27:72]
  wire  _T_687 = |alignicaf; // @[ifu_aln_ctl.scala 432:74]
  wire  _T_690 = first4B & _T_687; // @[Mux.scala 27:72]
  wire  _T_691 = first2B & alignicaf[0]; // @[Mux.scala 27:72]
  wire  _T_696 = first4B & _T_534; // @[ifu_aln_ctl.scala 434:54]
  wire  _T_698 = _T_696 & f0val[0]; // @[ifu_aln_ctl.scala 434:66]
  wire  _T_700 = ~alignicaf[0]; // @[ifu_aln_ctl.scala 434:79]
  wire  _T_701 = _T_698 & _T_700; // @[ifu_aln_ctl.scala 434:77]
  wire  _T_703 = ~aligndbecc[0]; // @[ifu_aln_ctl.scala 434:95]
  wire  _T_704 = _T_701 & _T_703; // @[ifu_aln_ctl.scala 434:93]
  wire [1:0] icaf_eff = alignicaf | aligndbecc; // @[ifu_aln_ctl.scala 436:28]
  wire  _T_708 = ~icaf_eff[0]; // @[ifu_aln_ctl.scala 438:53]
  wire  _T_709 = first4B & _T_708; // @[ifu_aln_ctl.scala 438:51]
  wire  _T_713 = |aligndbecc; // @[ifu_aln_ctl.scala 440:74]
  wire  _T_716 = first4B & _T_713; // @[Mux.scala 27:72]
  wire  _T_717 = first2B & aligndbecc[0]; // @[Mux.scala 27:72]
  wire [31:0] _T_726 = _T_682 ? aligndata : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_727 = _T_683 ? decompressed_io_dout : 32'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_732 = firstpc[8:1] ^ firstpc[16:9]; // @[lib.scala 51:47]
  wire [7:0] firstpc_hash = _T_732 ^ firstpc[24:17]; // @[lib.scala 51:85]
  wire [7:0] _T_736 = secondpc[8:1] ^ secondpc[16:9]; // @[lib.scala 51:47]
  wire [7:0] secondpc_hash = _T_736 ^ secondpc[24:17]; // @[lib.scala 51:85]
  wire [4:0] _T_742 = firstpc[13:9] ^ firstpc[18:14]; // @[lib.scala 42:111]
  wire [4:0] firstbrtag_hash = _T_742 ^ firstpc[23:19]; // @[lib.scala 42:111]
  wire [4:0] _T_748 = secondpc[13:9] ^ secondpc[18:14]; // @[lib.scala 42:111]
  wire [4:0] secondbrtag_hash = _T_748 ^ secondpc[23:19]; // @[lib.scala 42:111]
  wire  _T_751 = first2B & alignbrend[0]; // @[ifu_aln_ctl.scala 462:48]
  wire  _T_753 = first4B & alignbrend[1]; // @[ifu_aln_ctl.scala 462:76]
  wire  _T_754 = _T_751 | _T_753; // @[ifu_aln_ctl.scala 462:65]
  wire  _T_758 = _T_682 & alignbrend[0]; // @[ifu_aln_ctl.scala 462:118]
  wire  _T_761 = first2B & alignpc4[0]; // @[ifu_aln_ctl.scala 464:31]
  wire  _T_763 = first4B & alignpc4[1]; // @[ifu_aln_ctl.scala 464:57]
  wire  _T_764 = _T_761 | _T_763; // @[ifu_aln_ctl.scala 464:46]
  wire  _T_766 = first2B & alignret[0]; // @[ifu_aln_ctl.scala 466:51]
  wire  _T_768 = first4B & alignret[1]; // @[ifu_aln_ctl.scala 466:77]
  wire  _T_771 = first2B | alignbrend[0]; // @[ifu_aln_ctl.scala 468:55]
  wire  _T_777 = first2B & alignhist1[0]; // @[ifu_aln_ctl.scala 470:56]
  wire  _T_779 = first4B & alignhist1[1]; // @[ifu_aln_ctl.scala 470:84]
  wire  _T_780 = _T_777 | _T_779; // @[ifu_aln_ctl.scala 470:73]
  wire  _T_782 = first2B & alignhist0[0]; // @[ifu_aln_ctl.scala 471:16]
  wire  _T_784 = first4B & alignhist0[1]; // @[ifu_aln_ctl.scala 471:44]
  wire  _T_785 = _T_782 | _T_784; // @[ifu_aln_ctl.scala 471:33]
  wire  _T_787 = first4B & _T_536; // @[ifu_aln_ctl.scala 473:30]
  wire  _T_802 = io_dec_aln_aln_ib_i0_brp_valid & _T_764; // @[ifu_aln_ctl.scala 482:79]
  wire  _T_803 = _T_802 & first2B; // @[ifu_aln_ctl.scala 482:93]
  wire  _T_804 = ~_T_764; // @[ifu_aln_ctl.scala 482:141]
  wire  _T_805 = io_dec_aln_aln_ib_i0_brp_valid & _T_804; // @[ifu_aln_ctl.scala 482:139]
  wire  _T_806 = _T_805 & first4B; // @[ifu_aln_ctl.scala 482:153]
  wire [31:0] _T_820 = first2B ? aligndata : 32'h0; // @[ifu_aln_ctl.scala 502:29]
  rvclkhdr rvclkhdr ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en)
  );
  ifu_compress_ctl decompressed ( // @[ifu_aln_ctl.scala 444:28]
    .io_din(decompressed_io_din),
    .io_dout(decompressed_io_dout)
  );
  assign io_dec_aln_aln_dec_ifu_i0_cinst = aligndata[15:0]; // @[ifu_aln_ctl.scala 423:35]
  assign io_dec_aln_aln_ib_ifu_i0_icaf = _T_690 | _T_691; // @[ifu_aln_ctl.scala 432:33]
  assign io_dec_aln_aln_ib_ifu_i0_icaf_type = _T_704 ? f1ictype : f0ictype; // @[ifu_aln_ctl.scala 434:38]
  assign io_dec_aln_aln_ib_ifu_i0_icaf_second = _T_709 & icaf_eff[1]; // @[ifu_aln_ctl.scala 438:40]
  assign io_dec_aln_aln_ib_ifu_i0_dbecc = _T_716 | _T_717; // @[ifu_aln_ctl.scala 440:34]
  assign io_dec_aln_aln_ib_ifu_i0_bp_index = _T_771 ? firstpc_hash : secondpc_hash; // @[ifu_aln_ctl.scala 484:39]
  assign io_dec_aln_aln_ib_ifu_i0_bp_fghr = _T_787 ? f1fghr : f0fghr; // @[ifu_aln_ctl.scala 485:38]
  assign io_dec_aln_aln_ib_ifu_i0_bp_btag = _T_771 ? firstbrtag_hash : secondbrtag_hash; // @[ifu_aln_ctl.scala 486:38]
  assign io_dec_aln_aln_ib_ifu_i0_valid = _T_682 | _T_683; // @[ifu_aln_ctl.scala 430:34]
  assign io_dec_aln_aln_ib_ifu_i0_instr = _T_726 | _T_727; // @[ifu_aln_ctl.scala 446:34]
  assign io_dec_aln_aln_ib_ifu_i0_pc = _T_528 | _T_529; // @[ifu_aln_ctl.scala 419:31]
  assign io_dec_aln_aln_ib_ifu_i0_pc4 = aligndata[1:0] == 2'h3; // @[ifu_aln_ctl.scala 421:32]
  assign io_dec_aln_aln_ib_i0_brp_valid = _T_754 | _T_758; // @[ifu_aln_ctl.scala 462:36]
  assign io_dec_aln_aln_ib_i0_brp_bits_toffset = _T_787 ? f1poffset : f0poffset; // @[ifu_aln_ctl.scala 474:43]
  assign io_dec_aln_aln_ib_i0_brp_bits_hist = {_T_780,_T_785}; // @[ifu_aln_ctl.scala 470:40]
  assign io_dec_aln_aln_ib_i0_brp_bits_br_error = _T_803 | _T_806; // @[ifu_aln_ctl.scala 482:44]
  assign io_dec_aln_aln_ib_i0_brp_bits_br_start_error = _T_682 & alignbrend[0]; // @[ifu_aln_ctl.scala 478:51]
  assign io_dec_aln_aln_ib_i0_brp_bits_bank = _T_771 ? firstpc[0] : secondpc[0]; // @[ifu_aln_ctl.scala 480:51]
  assign io_dec_aln_aln_ib_i0_brp_bits_prett = _T_787 ? f1prett : f0prett; // @[ifu_aln_ctl.scala 476:41]
  assign io_dec_aln_aln_ib_i0_brp_bits_way = _T_771 ? alignway[0] : alignway[1]; // @[ifu_aln_ctl.scala 468:39]
  assign io_dec_aln_aln_ib_i0_brp_bits_ret = _T_766 | _T_768; // @[ifu_aln_ctl.scala 466:39]
  assign io_dec_aln_ifu_pmu_instr_aligned = io_dec_i0_decode_d & _T_821; // @[ifu_aln_ctl.scala 506:36]
  assign io_ifu_fb_consume1 = _T_350 & _T_1; // @[ifu_aln_ctl.scala 332:22]
  assign io_ifu_fb_consume2 = _T_353 & _T_1; // @[ifu_aln_ctl.scala 333:22]
  assign rvclkhdr_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_io_en = qwen[2]; // @[lib.scala 412:17]
  assign rvclkhdr_1_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_1_io_en = qwen[1]; // @[lib.scala 412:17]
  assign rvclkhdr_2_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_2_io_en = qwen[0]; // @[lib.scala 412:17]
  assign rvclkhdr_3_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_3_io_en = qwen[2]; // @[lib.scala 412:17]
  assign rvclkhdr_4_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_4_io_en = qwen[1]; // @[lib.scala 412:17]
  assign rvclkhdr_5_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_5_io_en = qwen[0]; // @[lib.scala 412:17]
  assign rvclkhdr_6_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_6_io_en = qwen[2]; // @[lib.scala 412:17]
  assign rvclkhdr_7_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_7_io_en = qwen[1]; // @[lib.scala 412:17]
  assign rvclkhdr_8_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_8_io_en = qwen[0]; // @[lib.scala 412:17]
  assign rvclkhdr_9_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_9_io_en = qwen[2]; // @[lib.scala 412:17]
  assign rvclkhdr_10_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_10_io_en = qwen[1]; // @[lib.scala 412:17]
  assign rvclkhdr_11_io_clk = clk; // @[lib.scala 411:18]
  assign rvclkhdr_11_io_en = qwen[0]; // @[lib.scala 412:17]
  assign decompressed_io_din = _T_820[15:0]; // @[ifu_aln_ctl.scala 502:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  error_stall = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wrptr = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  rdptr = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  q2off = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  q1off = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  q0off = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  f0val = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  q1 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  q0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  q2 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  f1val = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  f2val = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  brdata2 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  brdata1 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  brdata0 = _RAND_14[15:0];
  _RAND_15 = {2{`RANDOM}};
  misc2 = _RAND_15[52:0];
  _RAND_16 = {2{`RANDOM}};
  misc1 = _RAND_16[52:0];
  _RAND_17 = {2{`RANDOM}};
  misc0 = _RAND_17[52:0];
  _RAND_18 = {1{`RANDOM}};
  q2pc = _RAND_18[30:0];
  _RAND_19 = {1{`RANDOM}};
  q1pc = _RAND_19[30:0];
  _RAND_20 = {1{`RANDOM}};
  q0pc = _RAND_20[30:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    error_stall = 1'h0;
  end
  if (reset) begin
    wrptr = 2'h0;
  end
  if (reset) begin
    rdptr = 2'h0;
  end
  if (reset) begin
    q2off = 1'h0;
  end
  if (reset) begin
    q1off = 1'h0;
  end
  if (reset) begin
    q0off = 1'h0;
  end
  if (reset) begin
    f0val = 2'h0;
  end
  if (reset) begin
    q1 = 32'h0;
  end
  if (reset) begin
    q0 = 32'h0;
  end
  if (reset) begin
    q2 = 32'h0;
  end
  if (reset) begin
    f1val = 2'h0;
  end
  if (reset) begin
    f2val = 2'h0;
  end
  if (reset) begin
    brdata2 = 16'h0;
  end
  if (reset) begin
    brdata1 = 16'h0;
  end
  if (reset) begin
    brdata0 = 16'h0;
  end
  if (reset) begin
    misc2 = 53'h0;
  end
  if (reset) begin
    misc1 = 53'h0;
  end
  if (reset) begin
    misc0 = 53'h0;
  end
  if (reset) begin
    q2pc = 31'h0;
  end
  if (reset) begin
    q1pc = 31'h0;
  end
  if (reset) begin
    q0pc = 31'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      error_stall <= 1'h0;
    end else if (_T_4) begin
      error_stall <= error_stall_in;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      wrptr <= 2'h0;
    end else begin
      wrptr <= _T_118 | _T_117;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      rdptr <= 2'h0;
    end else begin
      rdptr <= _T_95 | _T_90;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      q2off <= 1'h0;
    end else begin
      q2off <= _T_142 | _T_141;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      q1off <= 1'h0;
    end else begin
      q1off <= _T_165 | _T_164;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      q0off <= 1'h0;
    end else begin
      q0off <= _T_188 | _T_187;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      f0val <= 2'h0;
    end else if (_T_13) begin
      f0val <= f0val_in;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      q1 <= 32'h0;
    end else if (qwen[1]) begin
      q1 <= io_ifu_fetch_data_f;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      q0 <= 32'h0;
    end else if (qwen[0]) begin
      q0 <= io_ifu_fetch_data_f;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      q2 <= 32'h0;
    end else if (qwen[2]) begin
      q2 <= io_ifu_fetch_data_f;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      f1val <= 2'h0;
    end else if (_T_10) begin
      f1val <= f1val_in;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      f2val <= 2'h0;
    end else if (_T_7) begin
      f2val <= f2val_in;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      brdata2 <= 16'h0;
    end else if (qwen[2]) begin
      brdata2 <= brdata_in;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      brdata1 <= 16'h0;
    end else if (qwen[1]) begin
      brdata1 <= brdata_in;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      brdata0 <= 16'h0;
    end else if (qwen[0]) begin
      brdata0 <= brdata_in;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      misc2 <= 53'h0;
    end else if (qwen[2]) begin
      misc2 <= misc_data_in;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      misc1 <= 53'h0;
    end else if (qwen[1]) begin
      misc1 <= misc_data_in;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      misc0 <= 53'h0;
    end else if (qwen[0]) begin
      misc0 <= misc_data_in;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      q2pc <= 31'h0;
    end else if (qwen[2]) begin
      q2pc <= io_ifu_fetch_pc;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      q1pc <= 31'h0;
    end else if (qwen[1]) begin
      q1pc <= io_ifu_fetch_pc;
    end
  end
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      q0pc <= 31'h0;
    end else if (qwen[0]) begin
      q0pc <= io_ifu_fetch_pc;
    end
  end
endmodule
module ifu_ifc_ctl(
  input         clock,
  input         reset,
  input         io_exu_flush_final,
  input  [30:0] io_exu_flush_path_final,
  input         io_free_l2clk,
  input         io_ic_hit_f,
  input         io_ifu_ic_mb_empty,
  input         io_ifu_fb_consume1,
  input         io_ifu_fb_consume2,
  input         io_ifu_bp_hit_taken_f,
  input  [30:0] io_ifu_bp_btb_target_f,
  input         io_ic_dma_active,
  input         io_ic_write_stall,
  input         io_dec_ifc_dec_tlu_flush_noredir_wb,
  input  [31:0] io_dec_ifc_dec_tlu_mrac_ff,
  output        io_dec_ifc_ifu_pmu_fetch_stall,
  input         io_dma_ifc_dma_iccm_stall_any,
  output [30:0] io_ifc_fetch_addr_f,
  output [30:0] io_ifc_fetch_addr_bf,
  output        io_ifc_fetch_req_f,
  output        io_ifc_fetch_uncacheable_bf,
  output        io_ifc_fetch_req_bf,
  output        io_ifc_fetch_req_bf_raw,
  output        io_ifc_iccm_access_bf,
  output        io_ifc_region_acc_fault_bf,
  output        io_ifc_dma_access_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg  dma_iccm_stall_any_f; // @[Reg.scala 27:20]
  wire  dma_stall = io_ic_dma_active | dma_iccm_stall_any_f; // @[ifu_ifc_ctl.scala 62:36]
  wire  _T_1 = io_dma_ifc_dma_iccm_stall_any ^ dma_iccm_stall_any_f; // @[lib.scala 475:21]
  wire  _T_2 = |_T_1; // @[lib.scala 475:29]
  wire  _T_56 = ~io_ic_hit_f; // @[ifu_ifc_ctl.scala 97:34]
  wire  _T_57 = io_ifc_fetch_req_f & _T_56; // @[ifu_ifc_ctl.scala 97:32]
  wire  _T_58 = ~io_exu_flush_final; // @[ifu_ifc_ctl.scala 97:49]
  wire  miss_f = _T_57 & _T_58; // @[ifu_ifc_ctl.scala 97:47]
  reg  miss_a; // @[Reg.scala 27:20]
  wire  _T_5 = miss_f ^ miss_a; // @[lib.scala 453:21]
  wire  _T_6 = |_T_5; // @[lib.scala 453:29]
  wire  _T_9 = ~io_ifc_fetch_req_f; // @[ifu_ifc_ctl.scala 67:53]
  wire  _T_11 = _T_9 | _T_56; // @[ifu_ifc_ctl.scala 67:73]
  wire  _T_12 = _T_58 & _T_11; // @[ifu_ifc_ctl.scala 67:50]
  wire  _T_14 = _T_58 & io_ifc_fetch_req_f; // @[ifu_ifc_ctl.scala 68:49]
  wire  _T_15 = _T_14 & io_ifu_bp_hit_taken_f; // @[ifu_ifc_ctl.scala 68:70]
  wire  _T_16 = _T_15 & io_ic_hit_f; // @[ifu_ifc_ctl.scala 68:94]
  wire  _T_19 = ~io_ifu_bp_hit_taken_f; // @[ifu_ifc_ctl.scala 69:73]
  wire  _T_20 = _T_14 & _T_19; // @[ifu_ifc_ctl.scala 69:71]
  wire  _T_21 = _T_20 & io_ic_hit_f; // @[ifu_ifc_ctl.scala 69:96]
  wire [30:0] _T_26 = io_exu_flush_final ? io_exu_flush_path_final : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_27 = _T_12 ? io_ifc_fetch_addr_f : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_28 = _T_16 ? io_ifu_bp_btb_target_f : 31'h0; // @[Mux.scala 27:72]
  wire [29:0] address_upper = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[ifu_ifc_ctl.scala 84:48]
  wire  _T_38 = address_upper[4] ^ io_ifc_fetch_addr_f[5]; // @[ifu_ifc_ctl.scala 85:63]
  wire  _T_39 = ~_T_38; // @[ifu_ifc_ctl.scala 85:24]
  wire  fetch_addr_next_0 = _T_39 & io_ifc_fetch_addr_f[0]; // @[ifu_ifc_ctl.scala 85:109]
  wire [30:0] fetch_addr_next = {address_upper,fetch_addr_next_0}; // @[Cat.scala 29:58]
  wire [30:0] _T_29 = _T_21 ? fetch_addr_next : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_30 = _T_26 | _T_27; // @[Mux.scala 27:72]
  wire [30:0] _T_31 = _T_30 | _T_28; // @[Mux.scala 27:72]
  reg [1:0] state; // @[Reg.scala 27:20]
  wire  idle = state == 2'h0; // @[ifu_ifc_ctl.scala 129:17]
  wire  _T_44 = io_ifu_fb_consume2 | io_ifu_fb_consume1; // @[ifu_ifc_ctl.scala 92:91]
  wire  _T_45 = ~_T_44; // @[ifu_ifc_ctl.scala 92:70]
  wire [3:0] _T_133 = io_exu_flush_final ? 4'h1 : 4'h0; // @[Mux.scala 27:72]
  wire  _T_93 = ~io_ifu_fb_consume2; // @[ifu_ifc_ctl.scala 115:38]
  wire  _T_94 = io_ifu_fb_consume1 & _T_93; // @[ifu_ifc_ctl.scala 115:36]
  wire  _T_96 = _T_9 | miss_f; // @[ifu_ifc_ctl.scala 115:81]
  wire  _T_97 = _T_94 & _T_96; // @[ifu_ifc_ctl.scala 115:58]
  wire  _T_98 = io_ifu_fb_consume2 & io_ifc_fetch_req_f; // @[ifu_ifc_ctl.scala 116:25]
  wire  fb_right = _T_97 | _T_98; // @[ifu_ifc_ctl.scala 115:92]
  wire  _T_110 = _T_58 & fb_right; // @[ifu_ifc_ctl.scala 123:16]
  reg [3:0] fb_write_f; // @[Reg.scala 27:20]
  wire [3:0] _T_113 = {1'h0,fb_write_f[3:1]}; // @[Cat.scala 29:58]
  wire [3:0] _T_134 = _T_110 ? _T_113 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_138 = _T_133 | _T_134; // @[Mux.scala 27:72]
  wire  fb_right2 = io_ifu_fb_consume2 & _T_96; // @[ifu_ifc_ctl.scala 118:36]
  wire  _T_115 = _T_58 & fb_right2; // @[ifu_ifc_ctl.scala 124:16]
  wire [3:0] _T_118 = {2'h0,fb_write_f[3:2]}; // @[Cat.scala 29:58]
  wire [3:0] _T_135 = _T_115 ? _T_118 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_139 = _T_138 | _T_135; // @[Mux.scala 27:72]
  wire  _T_103 = io_ifu_fb_consume1 | io_ifu_fb_consume2; // @[ifu_ifc_ctl.scala 119:56]
  wire  _T_104 = ~_T_103; // @[ifu_ifc_ctl.scala 119:35]
  wire  _T_105 = io_ifc_fetch_req_f & _T_104; // @[ifu_ifc_ctl.scala 119:33]
  wire  _T_106 = ~miss_f; // @[ifu_ifc_ctl.scala 119:80]
  wire  fb_left = _T_105 & _T_106; // @[ifu_ifc_ctl.scala 119:78]
  wire  _T_120 = _T_58 & fb_left; // @[ifu_ifc_ctl.scala 125:16]
  wire [3:0] _T_123 = {fb_write_f[2:0],1'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_136 = _T_120 ? _T_123 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_140 = _T_139 | _T_136; // @[Mux.scala 27:72]
  wire  _T_125 = ~fb_right; // @[ifu_ifc_ctl.scala 126:18]
  wire  _T_126 = _T_58 & _T_125; // @[ifu_ifc_ctl.scala 126:16]
  wire  _T_127 = ~fb_right2; // @[ifu_ifc_ctl.scala 126:30]
  wire  _T_128 = _T_126 & _T_127; // @[ifu_ifc_ctl.scala 126:28]
  wire  _T_129 = ~fb_left; // @[ifu_ifc_ctl.scala 126:43]
  wire  _T_130 = _T_128 & _T_129; // @[ifu_ifc_ctl.scala 126:41]
  wire [3:0] _T_137 = _T_130 ? fb_write_f : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] fb_write_ns = _T_140 | _T_137; // @[Mux.scala 27:72]
  wire  fb_full_f_ns = fb_write_ns[3]; // @[ifu_ifc_ctl.scala 132:30]
  wire  _T_46 = fb_full_f_ns & _T_45; // @[ifu_ifc_ctl.scala 92:68]
  wire  _T_47 = ~_T_46; // @[ifu_ifc_ctl.scala 92:53]
  wire  _T_48 = io_ifc_fetch_req_bf_raw & _T_47; // @[ifu_ifc_ctl.scala 92:51]
  wire  _T_49 = ~dma_stall; // @[ifu_ifc_ctl.scala 93:5]
  wire  _T_50 = _T_48 & _T_49; // @[ifu_ifc_ctl.scala 92:114]
  wire  _T_51 = ~io_ic_write_stall; // @[ifu_ifc_ctl.scala 93:18]
  wire  _T_52 = _T_50 & _T_51; // @[ifu_ifc_ctl.scala 93:16]
  wire  _T_53 = ~io_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu_ifc_ctl.scala 93:39]
  wire  fetch_bf_en = io_exu_flush_final | io_ifc_fetch_req_f; // @[ifu_ifc_ctl.scala 95:37]
  wire  _T_60 = io_ifu_ic_mb_empty | io_exu_flush_final; // @[ifu_ifc_ctl.scala 99:39]
  wire  _T_62 = _T_60 & _T_49; // @[ifu_ifc_ctl.scala 99:61]
  wire  _T_64 = _T_62 & _T_106; // @[ifu_ifc_ctl.scala 99:74]
  wire  _T_65 = ~miss_a; // @[ifu_ifc_ctl.scala 99:86]
  wire  mb_empty_mod = _T_64 & _T_65; // @[ifu_ifc_ctl.scala 99:84]
  wire  goto_idle = io_exu_flush_final & io_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu_ifc_ctl.scala 101:35]
  wire  _T_69 = io_exu_flush_final & _T_53; // @[ifu_ifc_ctl.scala 103:36]
  wire  leave_idle = _T_69 & idle; // @[ifu_ifc_ctl.scala 103:75]
  wire  _T_72 = ~state[1]; // @[ifu_ifc_ctl.scala 105:23]
  wire  _T_74 = _T_72 & state[0]; // @[ifu_ifc_ctl.scala 105:33]
  wire  _T_75 = _T_74 & miss_f; // @[ifu_ifc_ctl.scala 105:44]
  wire  _T_76 = ~goto_idle; // @[ifu_ifc_ctl.scala 105:55]
  wire  _T_77 = _T_75 & _T_76; // @[ifu_ifc_ctl.scala 105:53]
  wire  _T_79 = ~mb_empty_mod; // @[ifu_ifc_ctl.scala 106:17]
  wire  _T_80 = state[1] & _T_79; // @[ifu_ifc_ctl.scala 106:15]
  wire  _T_82 = _T_80 & _T_76; // @[ifu_ifc_ctl.scala 106:31]
  wire  next_state_1 = _T_77 | _T_82; // @[ifu_ifc_ctl.scala 105:67]
  wire  _T_84 = _T_76 & leave_idle; // @[ifu_ifc_ctl.scala 108:34]
  wire  _T_87 = state[0] & _T_76; // @[ifu_ifc_ctl.scala 108:60]
  wire  next_state_0 = _T_84 | _T_87; // @[ifu_ifc_ctl.scala 108:48]
  wire [1:0] _T_88 = {next_state_1,next_state_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_90 = _T_88 ^ state; // @[lib.scala 453:21]
  wire  _T_91 = |_T_90; // @[lib.scala 453:29]
  wire  wfm = state == 2'h3; // @[ifu_ifc_ctl.scala 130:16]
  reg  fb_full_f; // @[Reg.scala 27:20]
  wire  _T_146 = fb_full_f_ns ^ fb_full_f; // @[lib.scala 453:21]
  wire  _T_147 = |_T_146; // @[lib.scala 453:29]
  wire [3:0] _T_150 = fb_write_ns ^ fb_write_f; // @[lib.scala 453:21]
  wire  _T_151 = |_T_150; // @[lib.scala 453:29]
  wire  _T_154 = _T_44 | io_exu_flush_final; // @[ifu_ifc_ctl.scala 137:61]
  wire  _T_155 = ~_T_154; // @[ifu_ifc_ctl.scala 137:19]
  wire  _T_156 = fb_full_f & _T_155; // @[ifu_ifc_ctl.scala 137:17]
  wire  _T_157 = _T_156 | dma_stall; // @[ifu_ifc_ctl.scala 137:84]
  wire  _T_158 = io_ifc_fetch_req_bf_raw & _T_157; // @[ifu_ifc_ctl.scala 136:68]
  wire [31:0] _T_160 = {io_ifc_fetch_addr_bf,1'h0}; // @[Cat.scala 29:58]
  wire  iccm_acc_in_region_bf = _T_160[31:28] == 4'he; // @[lib.scala 84:47]
  wire  iccm_acc_in_range_bf = _T_160[31:16] == 16'hee00; // @[lib.scala 87:29]
  wire  _T_163 = ~io_ifc_iccm_access_bf; // @[ifu_ifc_ctl.scala 143:30]
  wire  _T_166 = fb_full_f & _T_45; // @[ifu_ifc_ctl.scala 144:16]
  wire  _T_167 = _T_163 | _T_166; // @[ifu_ifc_ctl.scala 143:53]
  wire  _T_168 = ~io_ifc_fetch_req_bf; // @[ifu_ifc_ctl.scala 145:13]
  wire  _T_169 = wfm & _T_168; // @[ifu_ifc_ctl.scala 145:11]
  wire  _T_170 = _T_167 | _T_169; // @[ifu_ifc_ctl.scala 144:62]
  wire  _T_171 = _T_170 | idle; // @[ifu_ifc_ctl.scala 145:35]
  wire  _T_173 = _T_171 & _T_58; // @[ifu_ifc_ctl.scala 145:44]
  wire  _T_175 = ~iccm_acc_in_range_bf; // @[ifu_ifc_ctl.scala 147:33]
  wire [4:0] _T_178 = {io_ifc_fetch_addr_bf[30:27],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_179 = io_dec_ifc_dec_tlu_mrac_ff >> _T_178; // @[ifu_ifc_ctl.scala 148:61]
  reg  _T_185; // @[Reg.scala 27:20]
  wire  _T_183 = io_ifc_fetch_req_bf ^ _T_185; // @[lib.scala 475:21]
  wire  _T_184 = |_T_183; // @[lib.scala 475:29]
  reg [30:0] _T_188; // @[Reg.scala 27:20]
  assign io_dec_ifc_ifu_pmu_fetch_stall = wfm | _T_158; // @[ifu_ifc_ctl.scala 136:34]
  assign io_ifc_fetch_addr_f = _T_188; // @[ifu_ifc_ctl.scala 152:23]
  assign io_ifc_fetch_addr_bf = _T_31 | _T_29; // @[ifu_ifc_ctl.scala 71:25]
  assign io_ifc_fetch_req_f = _T_185; // @[ifu_ifc_ctl.scala 150:22]
  assign io_ifc_fetch_uncacheable_bf = ~_T_179[0]; // @[ifu_ifc_ctl.scala 148:31]
  assign io_ifc_fetch_req_bf = _T_52 & _T_53; // @[ifu_ifc_ctl.scala 92:23]
  assign io_ifc_fetch_req_bf_raw = ~idle; // @[ifu_ifc_ctl.scala 90:27]
  assign io_ifc_iccm_access_bf = _T_160[31:16] == 16'hee00; // @[ifu_ifc_ctl.scala 142:25]
  assign io_ifc_region_acc_fault_bf = _T_175 & iccm_acc_in_region_bf; // @[ifu_ifc_ctl.scala 147:30]
  assign io_ifc_dma_access_ok = _T_173 | dma_iccm_stall_any_f; // @[ifu_ifc_ctl.scala 143:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dma_iccm_stall_any_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  miss_a = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  fb_write_f = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  fb_full_f = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_185 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_188 = _RAND_6[30:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    dma_iccm_stall_any_f = 1'h0;
  end
  if (reset) begin
    miss_a = 1'h0;
  end
  if (reset) begin
    state = 2'h0;
  end
  if (reset) begin
    fb_write_f = 4'h0;
  end
  if (reset) begin
    fb_full_f = 1'h0;
  end
  if (reset) begin
    _T_185 = 1'h0;
  end
  if (reset) begin
    _T_188 = 31'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      dma_iccm_stall_any_f <= 1'h0;
    end else if (_T_2) begin
      dma_iccm_stall_any_f <= io_dma_ifc_dma_iccm_stall_any;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      miss_a <= 1'h0;
    end else if (_T_6) begin
      miss_a <= miss_f;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_91) begin
      state <= _T_88;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      fb_write_f <= 4'h0;
    end else if (_T_151) begin
      fb_write_f <= fb_write_ns;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      fb_full_f <= 1'h0;
    end else if (_T_147) begin
      fb_full_f <= fb_full_f_ns;
    end
  end
  always @(posedge io_free_l2clk or posedge reset) begin
    if (reset) begin
      _T_185 <= 1'h0;
    end else if (_T_184) begin
      _T_185 <= io_ifc_fetch_req_bf;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_188 <= 31'h0;
    end else if (fetch_bf_en) begin
      _T_188 <= io_ifc_fetch_addr_bf;
    end
  end
endmodule
module ifu(
  input         clock,
  input         reset,
  output [8:0]  io_ifu_i0_fa_index,
  input         io_dec_i0_decode_d,
  input  [8:0]  io_dec_fa_error_index,
  input         io_exu_flush_final,
  input  [30:0] io_exu_flush_path_final,
  input         io_free_l2clk,
  input         io_active_clk,
  output [15:0] io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf,
  output [1:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_second,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc,
  output [7:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index,
  output [7:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr,
  output [4:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid,
  output [31:0] io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr,
  output [30:0] io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_valid,
  output [11:0] io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset,
  output [1:0]  io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_bank,
  output [30:0] io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret,
  output        io_ifu_dec_dec_aln_ifu_pmu_instr_aligned,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb,
  input  [70:0] io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_trxn,
  output        io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start,
  output        io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err,
  output [70:0] io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data,
  output        io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid,
  output        io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle,
  input         io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb,
  input  [31:0] io_ifu_dec_dec_ifc_dec_tlu_mrac_ff,
  output        io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid,
  input  [1:0]  io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle,
  input         io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb,
  input         io_ifu_dec_dec_bp_dec_tlu_bpred_disable,
  input  [7:0]  io_exu_ifu_exu_bp_exu_i0_br_index_r,
  input  [7:0]  io_exu_ifu_exu_bp_exu_i0_br_fghr_r,
  input         io_exu_ifu_exu_bp_exu_i0_br_way_r,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_valid,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_misp,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_ataken,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_boffset,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pc4,
  input  [1:0]  io_exu_ifu_exu_bp_exu_mp_pkt_bits_hist,
  input  [11:0] io_exu_ifu_exu_bp_exu_mp_pkt_bits_toffset,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_br_error,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_br_start_error,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pcall,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pja,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_way,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pret,
  input  [30:0] io_exu_ifu_exu_bp_exu_mp_pkt_bits_prett,
  input  [7:0]  io_exu_ifu_exu_bp_exu_mp_eghr,
  input  [7:0]  io_exu_ifu_exu_bp_exu_mp_fghr,
  input  [7:0]  io_exu_ifu_exu_bp_exu_mp_index,
  input  [4:0]  io_exu_ifu_exu_bp_exu_mp_btag,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [2:0]  io_iccm_wr_size,
  output [77:0] io_iccm_wr_data,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_tag_valid,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [9:0]  io_ic_debug_addr,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ic_tag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_ifu_aw_ready,
  output        io_ifu_aw_valid,
  output [2:0]  io_ifu_aw_bits_id,
  output [31:0] io_ifu_aw_bits_addr,
  output [3:0]  io_ifu_aw_bits_region,
  output [7:0]  io_ifu_aw_bits_len,
  output [2:0]  io_ifu_aw_bits_size,
  output [1:0]  io_ifu_aw_bits_burst,
  output        io_ifu_aw_bits_lock,
  output [3:0]  io_ifu_aw_bits_cache,
  output [2:0]  io_ifu_aw_bits_prot,
  output [3:0]  io_ifu_aw_bits_qos,
  input         io_ifu_w_ready,
  output        io_ifu_w_valid,
  output [63:0] io_ifu_w_bits_data,
  output [7:0]  io_ifu_w_bits_strb,
  output        io_ifu_w_bits_last,
  output        io_ifu_b_ready,
  input         io_ifu_b_valid,
  input  [1:0]  io_ifu_b_bits_resp,
  input  [2:0]  io_ifu_b_bits_id,
  input         io_ifu_ar_ready,
  output        io_ifu_ar_valid,
  output [2:0]  io_ifu_ar_bits_id,
  output [31:0] io_ifu_ar_bits_addr,
  output [3:0]  io_ifu_ar_bits_region,
  output [7:0]  io_ifu_ar_bits_len,
  output [2:0]  io_ifu_ar_bits_size,
  output [1:0]  io_ifu_ar_bits_burst,
  output        io_ifu_ar_bits_lock,
  output [3:0]  io_ifu_ar_bits_cache,
  output [2:0]  io_ifu_ar_bits_prot,
  output [3:0]  io_ifu_ar_bits_qos,
  output        io_ifu_r_ready,
  input         io_ifu_r_valid,
  input  [2:0]  io_ifu_r_bits_id,
  input  [63:0] io_ifu_r_bits_data,
  input  [1:0]  io_ifu_r_bits_resp,
  input         io_ifu_r_bits_last,
  input         io_ifu_bus_clk_en,
  input         io_ifu_dma_dma_ifc_dma_iccm_stall_any,
  input         io_ifu_dma_dma_mem_ctl_dma_iccm_req,
  input  [31:0] io_ifu_dma_dma_mem_ctl_dma_mem_addr,
  input  [2:0]  io_ifu_dma_dma_mem_ctl_dma_mem_sz,
  input         io_ifu_dma_dma_mem_ctl_dma_mem_write,
  input  [63:0] io_ifu_dma_dma_mem_ctl_dma_mem_wdata,
  input  [2:0]  io_ifu_dma_dma_mem_ctl_dma_mem_tag,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output        io_iccm_dma_sb_error,
  input         io_dec_tlu_flush_lower_wb,
  input         io_scan_mode
);
  wire  mem_ctl_clock; // @[ifu.scala 39:23]
  wire  mem_ctl_reset; // @[ifu.scala 39:23]
  wire  mem_ctl_io_free_l2clk; // @[ifu.scala 39:23]
  wire  mem_ctl_io_active_clk; // @[ifu.scala 39:23]
  wire  mem_ctl_io_exu_flush_final; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_fence_i_wb; // @[ifu.scala 39:23]
  wire [70:0] mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[ifu.scala 39:23]
  wire [16:0] mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_miss; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_hit; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_error; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_busy; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_trxn; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err; // @[ifu.scala 39:23]
  wire [70:0] mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_miss_state_idle; // @[ifu.scala 39:23]
  wire [30:0] mem_ctl_io_ifc_fetch_addr_bf; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifc_fetch_uncacheable_bf; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifc_fetch_req_bf; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifc_fetch_req_bf_raw; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifc_iccm_access_bf; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifc_region_acc_fault_bf; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifc_dma_access_ok; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifu_bp_inst_mask_f; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifu_axi_ar_ready; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifu_axi_ar_valid; // @[ifu.scala 39:23]
  wire [2:0] mem_ctl_io_ifu_axi_ar_bits_id; // @[ifu.scala 39:23]
  wire [31:0] mem_ctl_io_ifu_axi_ar_bits_addr; // @[ifu.scala 39:23]
  wire [3:0] mem_ctl_io_ifu_axi_ar_bits_region; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifu_axi_r_ready; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifu_axi_r_valid; // @[ifu.scala 39:23]
  wire [2:0] mem_ctl_io_ifu_axi_r_bits_id; // @[ifu.scala 39:23]
  wire [63:0] mem_ctl_io_ifu_axi_r_bits_data; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_ifu_axi_r_bits_resp; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifu_bus_clk_en; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dma_mem_ctl_dma_iccm_req; // @[ifu.scala 39:23]
  wire [31:0] mem_ctl_io_dma_mem_ctl_dma_mem_addr; // @[ifu.scala 39:23]
  wire [2:0] mem_ctl_io_dma_mem_ctl_dma_mem_sz; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dma_mem_ctl_dma_mem_write; // @[ifu.scala 39:23]
  wire [63:0] mem_ctl_io_dma_mem_ctl_dma_mem_wdata; // @[ifu.scala 39:23]
  wire [2:0] mem_ctl_io_dma_mem_ctl_dma_mem_tag; // @[ifu.scala 39:23]
  wire [14:0] mem_ctl_io_iccm_rw_addr; // @[ifu.scala 39:23]
  wire  mem_ctl_io_iccm_buf_correct_ecc; // @[ifu.scala 39:23]
  wire  mem_ctl_io_iccm_correction_state; // @[ifu.scala 39:23]
  wire  mem_ctl_io_iccm_wren; // @[ifu.scala 39:23]
  wire  mem_ctl_io_iccm_rden; // @[ifu.scala 39:23]
  wire [2:0] mem_ctl_io_iccm_wr_size; // @[ifu.scala 39:23]
  wire [77:0] mem_ctl_io_iccm_wr_data; // @[ifu.scala 39:23]
  wire [63:0] mem_ctl_io_iccm_rd_data; // @[ifu.scala 39:23]
  wire [77:0] mem_ctl_io_iccm_rd_data_ecc; // @[ifu.scala 39:23]
  wire [30:0] mem_ctl_io_ic_rw_addr; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_ic_tag_valid; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_ic_wr_en; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ic_rd_en; // @[ifu.scala 39:23]
  wire [70:0] mem_ctl_io_ic_wr_data_0; // @[ifu.scala 39:23]
  wire [70:0] mem_ctl_io_ic_wr_data_1; // @[ifu.scala 39:23]
  wire [70:0] mem_ctl_io_ic_debug_wr_data; // @[ifu.scala 39:23]
  wire [9:0] mem_ctl_io_ic_debug_addr; // @[ifu.scala 39:23]
  wire [63:0] mem_ctl_io_ic_rd_data; // @[ifu.scala 39:23]
  wire [70:0] mem_ctl_io_ic_debug_rd_data; // @[ifu.scala 39:23]
  wire [25:0] mem_ctl_io_ic_tag_debug_rd_data; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_ic_eccerr; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_ic_rd_hit; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ic_tag_perr; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ic_debug_rd_en; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ic_debug_wr_en; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ic_debug_tag_array; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_ic_debug_way; // @[ifu.scala 39:23]
  wire [63:0] mem_ctl_io_ic_premux_data; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ic_sel_premux_data; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_ifu_fetch_val; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifu_ic_mb_empty; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ic_dma_active; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ic_write_stall; // @[ifu.scala 39:23]
  wire  mem_ctl_io_iccm_dma_ecc_error; // @[ifu.scala 39:23]
  wire  mem_ctl_io_iccm_dma_rvalid; // @[ifu.scala 39:23]
  wire [63:0] mem_ctl_io_iccm_dma_rdata; // @[ifu.scala 39:23]
  wire [2:0] mem_ctl_io_iccm_dma_rtag; // @[ifu.scala 39:23]
  wire  mem_ctl_io_iccm_ready; // @[ifu.scala 39:23]
  wire  mem_ctl_io_dec_tlu_flush_lower_wb; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_iccm_rd_ecc_double_err; // @[ifu.scala 39:23]
  wire  mem_ctl_io_iccm_dma_sb_error; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ic_hit_f; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_ic_access_fault_f; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_ic_access_fault_type_f; // @[ifu.scala 39:23]
  wire  mem_ctl_io_ifu_async_error_start; // @[ifu.scala 39:23]
  wire [1:0] mem_ctl_io_ic_fetch_val_f; // @[ifu.scala 39:23]
  wire [31:0] mem_ctl_io_ic_data_f; // @[ifu.scala 39:23]
  wire  bp_ctl_clock; // @[ifu.scala 40:22]
  wire  bp_ctl_reset; // @[ifu.scala 40:22]
  wire  bp_ctl_io_ic_hit_f; // @[ifu.scala 40:22]
  wire  bp_ctl_io_exu_flush_final; // @[ifu.scala 40:22]
  wire [30:0] bp_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 40:22]
  wire  bp_ctl_io_ifc_fetch_req_f; // @[ifu.scala 40:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_valid; // @[ifu.scala 40:22]
  wire [1:0] bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_hist; // @[ifu.scala 40:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu.scala 40:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[ifu.scala 40:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu.scala 40:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu.scala 40:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_flush_leak_one_wb; // @[ifu.scala 40:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_bpred_disable; // @[ifu.scala 40:22]
  wire  bp_ctl_io_dec_tlu_flush_lower_wb; // @[ifu.scala 40:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_i0_br_index_r; // @[ifu.scala 40:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_i0_br_fghr_r; // @[ifu.scala 40:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_valid; // @[ifu.scala 40:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_misp; // @[ifu.scala 40:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu.scala 40:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu.scala 40:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pc4; // @[ifu.scala 40:22]
  wire [1:0] bp_ctl_io_exu_bp_exu_mp_pkt_bits_hist; // @[ifu.scala 40:22]
  wire [11:0] bp_ctl_io_exu_bp_exu_mp_pkt_bits_toffset; // @[ifu.scala 40:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu.scala 40:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu.scala 40:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_way; // @[ifu.scala 40:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pret; // @[ifu.scala 40:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_mp_eghr; // @[ifu.scala 40:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_mp_fghr; // @[ifu.scala 40:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_mp_index; // @[ifu.scala 40:22]
  wire [4:0] bp_ctl_io_exu_bp_exu_mp_btag; // @[ifu.scala 40:22]
  wire  bp_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 40:22]
  wire [30:0] bp_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 40:22]
  wire  bp_ctl_io_ifu_bp_inst_mask_f; // @[ifu.scala 40:22]
  wire [7:0] bp_ctl_io_ifu_bp_fghr_f; // @[ifu.scala 40:22]
  wire [1:0] bp_ctl_io_ifu_bp_way_f; // @[ifu.scala 40:22]
  wire [1:0] bp_ctl_io_ifu_bp_ret_f; // @[ifu.scala 40:22]
  wire [1:0] bp_ctl_io_ifu_bp_hist1_f; // @[ifu.scala 40:22]
  wire [1:0] bp_ctl_io_ifu_bp_hist0_f; // @[ifu.scala 40:22]
  wire [1:0] bp_ctl_io_ifu_bp_pc4_f; // @[ifu.scala 40:22]
  wire [1:0] bp_ctl_io_ifu_bp_valid_f; // @[ifu.scala 40:22]
  wire [11:0] bp_ctl_io_ifu_bp_poffset_f; // @[ifu.scala 40:22]
  wire  aln_ctl_clk; // @[ifu.scala 41:23]
  wire  aln_ctl_reset; // @[ifu.scala 41:23]
  wire  aln_ctl_io_active_clk; // @[ifu.scala 41:23]
  wire  aln_ctl_io_ifu_async_error_start; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_iccm_rd_ecc_double_err; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_ic_access_fault_f; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_ic_access_fault_type_f; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_i0_decode_d; // @[ifu.scala 41:23]
  wire [15:0] aln_ctl_io_dec_aln_aln_dec_ifu_i0_cinst; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_type; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_second; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_dbecc; // @[ifu.scala 41:23]
  wire [7:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_index; // @[ifu.scala 41:23]
  wire [7:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_fghr; // @[ifu.scala 41:23]
  wire [4:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_btag; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_valid; // @[ifu.scala 41:23]
  wire [31:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_instr; // @[ifu.scala 41:23]
  wire [30:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc4; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_valid; // @[ifu.scala 41:23]
  wire [11:0] aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_toffset; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_hist; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_error; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_start_error; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_bank; // @[ifu.scala 41:23]
  wire [30:0] aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_prett; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_way; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_ret; // @[ifu.scala 41:23]
  wire  aln_ctl_io_dec_aln_ifu_pmu_instr_aligned; // @[ifu.scala 41:23]
  wire [7:0] aln_ctl_io_ifu_bp_fghr_f; // @[ifu.scala 41:23]
  wire [30:0] aln_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 41:23]
  wire [11:0] aln_ctl_io_ifu_bp_poffset_f; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_ifu_bp_hist0_f; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_ifu_bp_hist1_f; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_ifu_bp_pc4_f; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_ifu_bp_way_f; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_ifu_bp_valid_f; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_ifu_bp_ret_f; // @[ifu.scala 41:23]
  wire  aln_ctl_io_exu_flush_final; // @[ifu.scala 41:23]
  wire [31:0] aln_ctl_io_ifu_fetch_data_f; // @[ifu.scala 41:23]
  wire [1:0] aln_ctl_io_ifu_fetch_val; // @[ifu.scala 41:23]
  wire [30:0] aln_ctl_io_ifu_fetch_pc; // @[ifu.scala 41:23]
  wire  aln_ctl_io_ifu_fb_consume1; // @[ifu.scala 41:23]
  wire  aln_ctl_io_ifu_fb_consume2; // @[ifu.scala 41:23]
  wire  ifc_ctl_clock; // @[ifu.scala 42:23]
  wire  ifc_ctl_reset; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_exu_flush_final; // @[ifu.scala 42:23]
  wire [30:0] ifc_ctl_io_exu_flush_path_final; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_free_l2clk; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ic_hit_f; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifu_ic_mb_empty; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifu_fb_consume1; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifu_fb_consume2; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 42:23]
  wire [30:0] ifc_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ic_dma_active; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ic_write_stall; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu.scala 42:23]
  wire [31:0] ifc_ctl_io_dec_ifc_dec_tlu_mrac_ff; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_dec_ifc_ifu_pmu_fetch_stall; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_dma_ifc_dma_iccm_stall_any; // @[ifu.scala 42:23]
  wire [30:0] ifc_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 42:23]
  wire [30:0] ifc_ctl_io_ifc_fetch_addr_bf; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifc_fetch_req_f; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifc_fetch_uncacheable_bf; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifc_fetch_req_bf; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifc_fetch_req_bf_raw; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifc_iccm_access_bf; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifc_region_acc_fault_bf; // @[ifu.scala 42:23]
  wire  ifc_ctl_io_ifc_dma_access_ok; // @[ifu.scala 42:23]
  ifu_mem_ctl mem_ctl ( // @[ifu.scala 39:23]
    .clock(mem_ctl_clock),
    .reset(mem_ctl_reset),
    .io_free_l2clk(mem_ctl_io_free_l2clk),
    .io_active_clk(mem_ctl_io_active_clk),
    .io_exu_flush_final(mem_ctl_io_exu_flush_final),
    .io_dec_mem_ctrl_dec_tlu_flush_err_wb(mem_ctl_io_dec_mem_ctrl_dec_tlu_flush_err_wb),
    .io_dec_mem_ctrl_dec_tlu_i0_commit_cmt(mem_ctl_io_dec_mem_ctrl_dec_tlu_i0_commit_cmt),
    .io_dec_mem_ctrl_dec_tlu_force_halt(mem_ctl_io_dec_mem_ctrl_dec_tlu_force_halt),
    .io_dec_mem_ctrl_dec_tlu_fence_i_wb(mem_ctl_io_dec_mem_ctrl_dec_tlu_fence_i_wb),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid),
    .io_dec_mem_ctrl_dec_tlu_core_ecc_disable(mem_ctl_io_dec_mem_ctrl_dec_tlu_core_ecc_disable),
    .io_dec_mem_ctrl_ifu_pmu_ic_miss(mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_miss),
    .io_dec_mem_ctrl_ifu_pmu_ic_hit(mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_hit),
    .io_dec_mem_ctrl_ifu_pmu_bus_error(mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_error),
    .io_dec_mem_ctrl_ifu_pmu_bus_busy(mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_busy),
    .io_dec_mem_ctrl_ifu_pmu_bus_trxn(mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_trxn),
    .io_dec_mem_ctrl_ifu_ic_error_start(mem_ctl_io_dec_mem_ctrl_ifu_ic_error_start),
    .io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err(mem_ctl_io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err),
    .io_dec_mem_ctrl_ifu_ic_debug_rd_data(mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data),
    .io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid(mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid),
    .io_dec_mem_ctrl_ifu_miss_state_idle(mem_ctl_io_dec_mem_ctrl_ifu_miss_state_idle),
    .io_ifc_fetch_addr_bf(mem_ctl_io_ifc_fetch_addr_bf),
    .io_ifc_fetch_uncacheable_bf(mem_ctl_io_ifc_fetch_uncacheable_bf),
    .io_ifc_fetch_req_bf(mem_ctl_io_ifc_fetch_req_bf),
    .io_ifc_fetch_req_bf_raw(mem_ctl_io_ifc_fetch_req_bf_raw),
    .io_ifc_iccm_access_bf(mem_ctl_io_ifc_iccm_access_bf),
    .io_ifc_region_acc_fault_bf(mem_ctl_io_ifc_region_acc_fault_bf),
    .io_ifc_dma_access_ok(mem_ctl_io_ifc_dma_access_ok),
    .io_ifu_bp_hit_taken_f(mem_ctl_io_ifu_bp_hit_taken_f),
    .io_ifu_bp_inst_mask_f(mem_ctl_io_ifu_bp_inst_mask_f),
    .io_ifu_axi_ar_ready(mem_ctl_io_ifu_axi_ar_ready),
    .io_ifu_axi_ar_valid(mem_ctl_io_ifu_axi_ar_valid),
    .io_ifu_axi_ar_bits_id(mem_ctl_io_ifu_axi_ar_bits_id),
    .io_ifu_axi_ar_bits_addr(mem_ctl_io_ifu_axi_ar_bits_addr),
    .io_ifu_axi_ar_bits_region(mem_ctl_io_ifu_axi_ar_bits_region),
    .io_ifu_axi_r_ready(mem_ctl_io_ifu_axi_r_ready),
    .io_ifu_axi_r_valid(mem_ctl_io_ifu_axi_r_valid),
    .io_ifu_axi_r_bits_id(mem_ctl_io_ifu_axi_r_bits_id),
    .io_ifu_axi_r_bits_data(mem_ctl_io_ifu_axi_r_bits_data),
    .io_ifu_axi_r_bits_resp(mem_ctl_io_ifu_axi_r_bits_resp),
    .io_ifu_bus_clk_en(mem_ctl_io_ifu_bus_clk_en),
    .io_dma_mem_ctl_dma_iccm_req(mem_ctl_io_dma_mem_ctl_dma_iccm_req),
    .io_dma_mem_ctl_dma_mem_addr(mem_ctl_io_dma_mem_ctl_dma_mem_addr),
    .io_dma_mem_ctl_dma_mem_sz(mem_ctl_io_dma_mem_ctl_dma_mem_sz),
    .io_dma_mem_ctl_dma_mem_write(mem_ctl_io_dma_mem_ctl_dma_mem_write),
    .io_dma_mem_ctl_dma_mem_wdata(mem_ctl_io_dma_mem_ctl_dma_mem_wdata),
    .io_dma_mem_ctl_dma_mem_tag(mem_ctl_io_dma_mem_ctl_dma_mem_tag),
    .io_iccm_rw_addr(mem_ctl_io_iccm_rw_addr),
    .io_iccm_buf_correct_ecc(mem_ctl_io_iccm_buf_correct_ecc),
    .io_iccm_correction_state(mem_ctl_io_iccm_correction_state),
    .io_iccm_wren(mem_ctl_io_iccm_wren),
    .io_iccm_rden(mem_ctl_io_iccm_rden),
    .io_iccm_wr_size(mem_ctl_io_iccm_wr_size),
    .io_iccm_wr_data(mem_ctl_io_iccm_wr_data),
    .io_iccm_rd_data(mem_ctl_io_iccm_rd_data),
    .io_iccm_rd_data_ecc(mem_ctl_io_iccm_rd_data_ecc),
    .io_ic_rw_addr(mem_ctl_io_ic_rw_addr),
    .io_ic_tag_valid(mem_ctl_io_ic_tag_valid),
    .io_ic_wr_en(mem_ctl_io_ic_wr_en),
    .io_ic_rd_en(mem_ctl_io_ic_rd_en),
    .io_ic_wr_data_0(mem_ctl_io_ic_wr_data_0),
    .io_ic_wr_data_1(mem_ctl_io_ic_wr_data_1),
    .io_ic_debug_wr_data(mem_ctl_io_ic_debug_wr_data),
    .io_ic_debug_addr(mem_ctl_io_ic_debug_addr),
    .io_ic_rd_data(mem_ctl_io_ic_rd_data),
    .io_ic_debug_rd_data(mem_ctl_io_ic_debug_rd_data),
    .io_ic_tag_debug_rd_data(mem_ctl_io_ic_tag_debug_rd_data),
    .io_ic_eccerr(mem_ctl_io_ic_eccerr),
    .io_ic_rd_hit(mem_ctl_io_ic_rd_hit),
    .io_ic_tag_perr(mem_ctl_io_ic_tag_perr),
    .io_ic_debug_rd_en(mem_ctl_io_ic_debug_rd_en),
    .io_ic_debug_wr_en(mem_ctl_io_ic_debug_wr_en),
    .io_ic_debug_tag_array(mem_ctl_io_ic_debug_tag_array),
    .io_ic_debug_way(mem_ctl_io_ic_debug_way),
    .io_ic_premux_data(mem_ctl_io_ic_premux_data),
    .io_ic_sel_premux_data(mem_ctl_io_ic_sel_premux_data),
    .io_ifu_fetch_val(mem_ctl_io_ifu_fetch_val),
    .io_ifu_ic_mb_empty(mem_ctl_io_ifu_ic_mb_empty),
    .io_ic_dma_active(mem_ctl_io_ic_dma_active),
    .io_ic_write_stall(mem_ctl_io_ic_write_stall),
    .io_iccm_dma_ecc_error(mem_ctl_io_iccm_dma_ecc_error),
    .io_iccm_dma_rvalid(mem_ctl_io_iccm_dma_rvalid),
    .io_iccm_dma_rdata(mem_ctl_io_iccm_dma_rdata),
    .io_iccm_dma_rtag(mem_ctl_io_iccm_dma_rtag),
    .io_iccm_ready(mem_ctl_io_iccm_ready),
    .io_dec_tlu_flush_lower_wb(mem_ctl_io_dec_tlu_flush_lower_wb),
    .io_iccm_rd_ecc_double_err(mem_ctl_io_iccm_rd_ecc_double_err),
    .io_iccm_dma_sb_error(mem_ctl_io_iccm_dma_sb_error),
    .io_ic_hit_f(mem_ctl_io_ic_hit_f),
    .io_ic_access_fault_f(mem_ctl_io_ic_access_fault_f),
    .io_ic_access_fault_type_f(mem_ctl_io_ic_access_fault_type_f),
    .io_ifu_async_error_start(mem_ctl_io_ifu_async_error_start),
    .io_ic_fetch_val_f(mem_ctl_io_ic_fetch_val_f),
    .io_ic_data_f(mem_ctl_io_ic_data_f)
  );
  ifu_bp_ctl bp_ctl ( // @[ifu.scala 40:22]
    .clock(bp_ctl_clock),
    .reset(bp_ctl_reset),
    .io_ic_hit_f(bp_ctl_io_ic_hit_f),
    .io_exu_flush_final(bp_ctl_io_exu_flush_final),
    .io_ifc_fetch_addr_f(bp_ctl_io_ifc_fetch_addr_f),
    .io_ifc_fetch_req_f(bp_ctl_io_ifc_fetch_req_f),
    .io_dec_bp_dec_tlu_br0_r_pkt_valid(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_valid),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_hist(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_hist),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_way(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_way),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_middle(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_middle),
    .io_dec_bp_dec_tlu_flush_leak_one_wb(bp_ctl_io_dec_bp_dec_tlu_flush_leak_one_wb),
    .io_dec_bp_dec_tlu_bpred_disable(bp_ctl_io_dec_bp_dec_tlu_bpred_disable),
    .io_dec_tlu_flush_lower_wb(bp_ctl_io_dec_tlu_flush_lower_wb),
    .io_exu_bp_exu_i0_br_index_r(bp_ctl_io_exu_bp_exu_i0_br_index_r),
    .io_exu_bp_exu_i0_br_fghr_r(bp_ctl_io_exu_bp_exu_i0_br_fghr_r),
    .io_exu_bp_exu_mp_pkt_valid(bp_ctl_io_exu_bp_exu_mp_pkt_valid),
    .io_exu_bp_exu_mp_pkt_bits_misp(bp_ctl_io_exu_bp_exu_mp_pkt_bits_misp),
    .io_exu_bp_exu_mp_pkt_bits_ataken(bp_ctl_io_exu_bp_exu_mp_pkt_bits_ataken),
    .io_exu_bp_exu_mp_pkt_bits_boffset(bp_ctl_io_exu_bp_exu_mp_pkt_bits_boffset),
    .io_exu_bp_exu_mp_pkt_bits_pc4(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pc4),
    .io_exu_bp_exu_mp_pkt_bits_hist(bp_ctl_io_exu_bp_exu_mp_pkt_bits_hist),
    .io_exu_bp_exu_mp_pkt_bits_toffset(bp_ctl_io_exu_bp_exu_mp_pkt_bits_toffset),
    .io_exu_bp_exu_mp_pkt_bits_pcall(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pcall),
    .io_exu_bp_exu_mp_pkt_bits_pja(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pja),
    .io_exu_bp_exu_mp_pkt_bits_way(bp_ctl_io_exu_bp_exu_mp_pkt_bits_way),
    .io_exu_bp_exu_mp_pkt_bits_pret(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pret),
    .io_exu_bp_exu_mp_eghr(bp_ctl_io_exu_bp_exu_mp_eghr),
    .io_exu_bp_exu_mp_fghr(bp_ctl_io_exu_bp_exu_mp_fghr),
    .io_exu_bp_exu_mp_index(bp_ctl_io_exu_bp_exu_mp_index),
    .io_exu_bp_exu_mp_btag(bp_ctl_io_exu_bp_exu_mp_btag),
    .io_ifu_bp_hit_taken_f(bp_ctl_io_ifu_bp_hit_taken_f),
    .io_ifu_bp_btb_target_f(bp_ctl_io_ifu_bp_btb_target_f),
    .io_ifu_bp_inst_mask_f(bp_ctl_io_ifu_bp_inst_mask_f),
    .io_ifu_bp_fghr_f(bp_ctl_io_ifu_bp_fghr_f),
    .io_ifu_bp_way_f(bp_ctl_io_ifu_bp_way_f),
    .io_ifu_bp_ret_f(bp_ctl_io_ifu_bp_ret_f),
    .io_ifu_bp_hist1_f(bp_ctl_io_ifu_bp_hist1_f),
    .io_ifu_bp_hist0_f(bp_ctl_io_ifu_bp_hist0_f),
    .io_ifu_bp_pc4_f(bp_ctl_io_ifu_bp_pc4_f),
    .io_ifu_bp_valid_f(bp_ctl_io_ifu_bp_valid_f),
    .io_ifu_bp_poffset_f(bp_ctl_io_ifu_bp_poffset_f)
  );
  ifu_aln_ctl aln_ctl ( // @[ifu.scala 41:23]
    .clk(aln_ctl_clk),
    .reset(aln_ctl_reset),
    .io_active_clk(aln_ctl_io_active_clk),
    .io_ifu_async_error_start(aln_ctl_io_ifu_async_error_start),
    .io_iccm_rd_ecc_double_err(aln_ctl_io_iccm_rd_ecc_double_err),
    .io_ic_access_fault_f(aln_ctl_io_ic_access_fault_f),
    .io_ic_access_fault_type_f(aln_ctl_io_ic_access_fault_type_f),
    .io_dec_i0_decode_d(aln_ctl_io_dec_i0_decode_d),
    .io_dec_aln_aln_dec_ifu_i0_cinst(aln_ctl_io_dec_aln_aln_dec_ifu_i0_cinst),
    .io_dec_aln_aln_ib_ifu_i0_icaf(aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf),
    .io_dec_aln_aln_ib_ifu_i0_icaf_type(aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_type),
    .io_dec_aln_aln_ib_ifu_i0_icaf_second(aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_second),
    .io_dec_aln_aln_ib_ifu_i0_dbecc(aln_ctl_io_dec_aln_aln_ib_ifu_i0_dbecc),
    .io_dec_aln_aln_ib_ifu_i0_bp_index(aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_index),
    .io_dec_aln_aln_ib_ifu_i0_bp_fghr(aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_fghr),
    .io_dec_aln_aln_ib_ifu_i0_bp_btag(aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_btag),
    .io_dec_aln_aln_ib_ifu_i0_valid(aln_ctl_io_dec_aln_aln_ib_ifu_i0_valid),
    .io_dec_aln_aln_ib_ifu_i0_instr(aln_ctl_io_dec_aln_aln_ib_ifu_i0_instr),
    .io_dec_aln_aln_ib_ifu_i0_pc(aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc),
    .io_dec_aln_aln_ib_ifu_i0_pc4(aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc4),
    .io_dec_aln_aln_ib_i0_brp_valid(aln_ctl_io_dec_aln_aln_ib_i0_brp_valid),
    .io_dec_aln_aln_ib_i0_brp_bits_toffset(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_toffset),
    .io_dec_aln_aln_ib_i0_brp_bits_hist(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_hist),
    .io_dec_aln_aln_ib_i0_brp_bits_br_error(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_error),
    .io_dec_aln_aln_ib_i0_brp_bits_br_start_error(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_start_error),
    .io_dec_aln_aln_ib_i0_brp_bits_bank(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_bank),
    .io_dec_aln_aln_ib_i0_brp_bits_prett(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_prett),
    .io_dec_aln_aln_ib_i0_brp_bits_way(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_way),
    .io_dec_aln_aln_ib_i0_brp_bits_ret(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_ret),
    .io_dec_aln_ifu_pmu_instr_aligned(aln_ctl_io_dec_aln_ifu_pmu_instr_aligned),
    .io_ifu_bp_fghr_f(aln_ctl_io_ifu_bp_fghr_f),
    .io_ifu_bp_btb_target_f(aln_ctl_io_ifu_bp_btb_target_f),
    .io_ifu_bp_poffset_f(aln_ctl_io_ifu_bp_poffset_f),
    .io_ifu_bp_hist0_f(aln_ctl_io_ifu_bp_hist0_f),
    .io_ifu_bp_hist1_f(aln_ctl_io_ifu_bp_hist1_f),
    .io_ifu_bp_pc4_f(aln_ctl_io_ifu_bp_pc4_f),
    .io_ifu_bp_way_f(aln_ctl_io_ifu_bp_way_f),
    .io_ifu_bp_valid_f(aln_ctl_io_ifu_bp_valid_f),
    .io_ifu_bp_ret_f(aln_ctl_io_ifu_bp_ret_f),
    .io_exu_flush_final(aln_ctl_io_exu_flush_final),
    .io_ifu_fetch_data_f(aln_ctl_io_ifu_fetch_data_f),
    .io_ifu_fetch_val(aln_ctl_io_ifu_fetch_val),
    .io_ifu_fetch_pc(aln_ctl_io_ifu_fetch_pc),
    .io_ifu_fb_consume1(aln_ctl_io_ifu_fb_consume1),
    .io_ifu_fb_consume2(aln_ctl_io_ifu_fb_consume2)
  );
  ifu_ifc_ctl ifc_ctl ( // @[ifu.scala 42:23]
    .clock(ifc_ctl_clock),
    .reset(ifc_ctl_reset),
    .io_exu_flush_final(ifc_ctl_io_exu_flush_final),
    .io_exu_flush_path_final(ifc_ctl_io_exu_flush_path_final),
    .io_free_l2clk(ifc_ctl_io_free_l2clk),
    .io_ic_hit_f(ifc_ctl_io_ic_hit_f),
    .io_ifu_ic_mb_empty(ifc_ctl_io_ifu_ic_mb_empty),
    .io_ifu_fb_consume1(ifc_ctl_io_ifu_fb_consume1),
    .io_ifu_fb_consume2(ifc_ctl_io_ifu_fb_consume2),
    .io_ifu_bp_hit_taken_f(ifc_ctl_io_ifu_bp_hit_taken_f),
    .io_ifu_bp_btb_target_f(ifc_ctl_io_ifu_bp_btb_target_f),
    .io_ic_dma_active(ifc_ctl_io_ic_dma_active),
    .io_ic_write_stall(ifc_ctl_io_ic_write_stall),
    .io_dec_ifc_dec_tlu_flush_noredir_wb(ifc_ctl_io_dec_ifc_dec_tlu_flush_noredir_wb),
    .io_dec_ifc_dec_tlu_mrac_ff(ifc_ctl_io_dec_ifc_dec_tlu_mrac_ff),
    .io_dec_ifc_ifu_pmu_fetch_stall(ifc_ctl_io_dec_ifc_ifu_pmu_fetch_stall),
    .io_dma_ifc_dma_iccm_stall_any(ifc_ctl_io_dma_ifc_dma_iccm_stall_any),
    .io_ifc_fetch_addr_f(ifc_ctl_io_ifc_fetch_addr_f),
    .io_ifc_fetch_addr_bf(ifc_ctl_io_ifc_fetch_addr_bf),
    .io_ifc_fetch_req_f(ifc_ctl_io_ifc_fetch_req_f),
    .io_ifc_fetch_uncacheable_bf(ifc_ctl_io_ifc_fetch_uncacheable_bf),
    .io_ifc_fetch_req_bf(ifc_ctl_io_ifc_fetch_req_bf),
    .io_ifc_fetch_req_bf_raw(ifc_ctl_io_ifc_fetch_req_bf_raw),
    .io_ifc_iccm_access_bf(ifc_ctl_io_ifc_iccm_access_bf),
    .io_ifc_region_acc_fault_bf(ifc_ctl_io_ifc_region_acc_fault_bf),
    .io_ifc_dma_access_ok(ifc_ctl_io_ifc_dma_access_ok)
  );
  assign io_ifu_i0_fa_index = 9'h0; // @[ifu.scala 85:56]
  assign io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst = aln_ctl_io_dec_aln_aln_dec_ifu_i0_cinst; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf = aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type = aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_type; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_second = aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_second; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc = aln_ctl_io_dec_aln_aln_ib_ifu_i0_dbecc; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index = aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_index; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr = aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_fghr; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag = aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_btag; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid = aln_ctl_io_dec_aln_aln_ib_ifu_i0_valid; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr = aln_ctl_io_dec_aln_aln_ib_ifu_i0_instr; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc = aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4 = aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc4; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_valid = aln_ctl_io_dec_aln_aln_ib_i0_brp_valid; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_toffset; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_hist; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_error; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_start_error; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_bank = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_bank; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_prett; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_way; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_ret; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_aln_ifu_pmu_instr_aligned = aln_ctl_io_dec_aln_ifu_pmu_instr_aligned; // @[ifu.scala 78:22]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss = mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_miss; // @[ifu.scala 117:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit = mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_hit; // @[ifu.scala 117:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error = mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_error; // @[ifu.scala 117:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy = mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_busy; // @[ifu.scala 117:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_trxn = mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_trxn; // @[ifu.scala 117:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start = mem_ctl_io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu.scala 117:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err = mem_ctl_io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err; // @[ifu.scala 117:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data = mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data; // @[ifu.scala 117:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid = mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid; // @[ifu.scala 117:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle = mem_ctl_io_dec_mem_ctrl_ifu_miss_state_idle; // @[ifu.scala 117:27]
  assign io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall = ifc_ctl_io_dec_ifc_ifu_pmu_fetch_stall; // @[ifu.scala 51:22]
  assign io_iccm_rw_addr = mem_ctl_io_iccm_rw_addr; // @[ifu.scala 131:19]
  assign io_iccm_buf_correct_ecc = mem_ctl_io_iccm_buf_correct_ecc; // @[ifu.scala 131:19]
  assign io_iccm_correction_state = mem_ctl_io_iccm_correction_state; // @[ifu.scala 131:19]
  assign io_iccm_wren = mem_ctl_io_iccm_wren; // @[ifu.scala 131:19]
  assign io_iccm_rden = mem_ctl_io_iccm_rden; // @[ifu.scala 131:19]
  assign io_iccm_wr_size = mem_ctl_io_iccm_wr_size; // @[ifu.scala 131:19]
  assign io_iccm_wr_data = mem_ctl_io_iccm_wr_data; // @[ifu.scala 131:19]
  assign io_ic_rw_addr = mem_ctl_io_ic_rw_addr; // @[ifu.scala 130:17]
  assign io_ic_tag_valid = mem_ctl_io_ic_tag_valid; // @[ifu.scala 130:17]
  assign io_ic_wr_en = mem_ctl_io_ic_wr_en; // @[ifu.scala 130:17]
  assign io_ic_rd_en = mem_ctl_io_ic_rd_en; // @[ifu.scala 130:17]
  assign io_ic_wr_data_0 = mem_ctl_io_ic_wr_data_0; // @[ifu.scala 130:17]
  assign io_ic_wr_data_1 = mem_ctl_io_ic_wr_data_1; // @[ifu.scala 130:17]
  assign io_ic_debug_wr_data = mem_ctl_io_ic_debug_wr_data; // @[ifu.scala 130:17]
  assign io_ic_debug_addr = mem_ctl_io_ic_debug_addr; // @[ifu.scala 130:17]
  assign io_ic_debug_rd_en = mem_ctl_io_ic_debug_rd_en; // @[ifu.scala 130:17]
  assign io_ic_debug_wr_en = mem_ctl_io_ic_debug_wr_en; // @[ifu.scala 130:17]
  assign io_ic_debug_tag_array = mem_ctl_io_ic_debug_tag_array; // @[ifu.scala 130:17]
  assign io_ic_debug_way = mem_ctl_io_ic_debug_way; // @[ifu.scala 130:17]
  assign io_ic_premux_data = mem_ctl_io_ic_premux_data; // @[ifu.scala 130:17]
  assign io_ic_sel_premux_data = mem_ctl_io_ic_sel_premux_data; // @[ifu.scala 130:17]
  assign io_ifu_aw_valid = 1'h0; // @[ifu.scala 127:22]
  assign io_ifu_aw_bits_id = 3'h0; // @[ifu.scala 127:22]
  assign io_ifu_aw_bits_addr = 32'h0; // @[ifu.scala 127:22]
  assign io_ifu_aw_bits_region = 4'h0; // @[ifu.scala 127:22]
  assign io_ifu_aw_bits_len = 8'h0; // @[ifu.scala 127:22]
  assign io_ifu_aw_bits_size = 3'h0; // @[ifu.scala 127:22]
  assign io_ifu_aw_bits_burst = 2'h0; // @[ifu.scala 127:22]
  assign io_ifu_aw_bits_lock = 1'h0; // @[ifu.scala 127:22]
  assign io_ifu_aw_bits_cache = 4'h0; // @[ifu.scala 127:22]
  assign io_ifu_aw_bits_prot = 3'h0; // @[ifu.scala 127:22]
  assign io_ifu_aw_bits_qos = 4'h0; // @[ifu.scala 127:22]
  assign io_ifu_w_valid = 1'h0; // @[ifu.scala 127:22]
  assign io_ifu_w_bits_data = 64'h0; // @[ifu.scala 127:22]
  assign io_ifu_w_bits_strb = 8'h0; // @[ifu.scala 127:22]
  assign io_ifu_w_bits_last = 1'h0; // @[ifu.scala 127:22]
  assign io_ifu_b_ready = 1'h0; // @[ifu.scala 127:22]
  assign io_ifu_ar_valid = mem_ctl_io_ifu_axi_ar_valid; // @[ifu.scala 127:22]
  assign io_ifu_ar_bits_id = mem_ctl_io_ifu_axi_ar_bits_id; // @[ifu.scala 127:22]
  assign io_ifu_ar_bits_addr = mem_ctl_io_ifu_axi_ar_bits_addr; // @[ifu.scala 127:22]
  assign io_ifu_ar_bits_region = mem_ctl_io_ifu_axi_ar_bits_region; // @[ifu.scala 127:22]
  assign io_ifu_ar_bits_len = 8'h0; // @[ifu.scala 127:22]
  assign io_ifu_ar_bits_size = 3'h3; // @[ifu.scala 127:22]
  assign io_ifu_ar_bits_burst = 2'h1; // @[ifu.scala 127:22]
  assign io_ifu_ar_bits_lock = 1'h0; // @[ifu.scala 127:22]
  assign io_ifu_ar_bits_cache = 4'hf; // @[ifu.scala 127:22]
  assign io_ifu_ar_bits_prot = 3'h5; // @[ifu.scala 127:22]
  assign io_ifu_ar_bits_qos = 4'h0; // @[ifu.scala 127:22]
  assign io_ifu_r_ready = 1'h1; // @[ifu.scala 127:22]
  assign io_iccm_dma_ecc_error = mem_ctl_io_iccm_dma_ecc_error; // @[ifu.scala 137:25]
  assign io_iccm_dma_rvalid = mem_ctl_io_iccm_dma_rvalid; // @[ifu.scala 138:22]
  assign io_iccm_dma_rdata = mem_ctl_io_iccm_dma_rdata; // @[ifu.scala 139:21]
  assign io_iccm_dma_rtag = mem_ctl_io_iccm_dma_rtag; // @[ifu.scala 140:20]
  assign io_iccm_ready = mem_ctl_io_iccm_ready; // @[ifu.scala 141:17]
  assign io_iccm_dma_sb_error = mem_ctl_io_iccm_dma_sb_error; // @[ifu.scala 142:24]
  assign mem_ctl_clock = clock;
  assign mem_ctl_reset = reset;
  assign mem_ctl_io_free_l2clk = io_free_l2clk; // @[ifu.scala 114:25]
  assign mem_ctl_io_active_clk = io_active_clk; // @[ifu.scala 115:25]
  assign mem_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 116:30]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_flush_err_wb = io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu.scala 117:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_i0_commit_cmt = io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu.scala 117:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_force_halt = io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu.scala 117:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_fence_i_wb = io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb; // @[ifu.scala 117:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[ifu.scala 117:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics; // @[ifu.scala 117:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[ifu.scala 117:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[ifu.scala 117:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_core_ecc_disable = io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[ifu.scala 117:27]
  assign mem_ctl_io_ifc_fetch_addr_bf = ifc_ctl_io_ifc_fetch_addr_bf; // @[ifu.scala 118:32]
  assign mem_ctl_io_ifc_fetch_uncacheable_bf = ifc_ctl_io_ifc_fetch_uncacheable_bf; // @[ifu.scala 119:39]
  assign mem_ctl_io_ifc_fetch_req_bf = ifc_ctl_io_ifc_fetch_req_bf; // @[ifu.scala 120:31]
  assign mem_ctl_io_ifc_fetch_req_bf_raw = ifc_ctl_io_ifc_fetch_req_bf_raw; // @[ifu.scala 121:35]
  assign mem_ctl_io_ifc_iccm_access_bf = ifc_ctl_io_ifc_iccm_access_bf; // @[ifu.scala 122:33]
  assign mem_ctl_io_ifc_region_acc_fault_bf = ifc_ctl_io_ifc_region_acc_fault_bf; // @[ifu.scala 123:38]
  assign mem_ctl_io_ifc_dma_access_ok = ifc_ctl_io_ifc_dma_access_ok; // @[ifu.scala 124:32]
  assign mem_ctl_io_ifu_bp_hit_taken_f = bp_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 125:33]
  assign mem_ctl_io_ifu_bp_inst_mask_f = bp_ctl_io_ifu_bp_inst_mask_f; // @[ifu.scala 126:33]
  assign mem_ctl_io_ifu_axi_ar_ready = io_ifu_ar_ready; // @[ifu.scala 127:22]
  assign mem_ctl_io_ifu_axi_r_valid = io_ifu_r_valid; // @[ifu.scala 127:22]
  assign mem_ctl_io_ifu_axi_r_bits_id = io_ifu_r_bits_id; // @[ifu.scala 127:22]
  assign mem_ctl_io_ifu_axi_r_bits_data = io_ifu_r_bits_data; // @[ifu.scala 127:22]
  assign mem_ctl_io_ifu_axi_r_bits_resp = io_ifu_r_bits_resp; // @[ifu.scala 127:22]
  assign mem_ctl_io_ifu_bus_clk_en = io_ifu_bus_clk_en; // @[ifu.scala 128:29]
  assign mem_ctl_io_dma_mem_ctl_dma_iccm_req = io_ifu_dma_dma_mem_ctl_dma_iccm_req; // @[ifu.scala 129:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_addr = io_ifu_dma_dma_mem_ctl_dma_mem_addr; // @[ifu.scala 129:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_sz = io_ifu_dma_dma_mem_ctl_dma_mem_sz; // @[ifu.scala 129:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_write = io_ifu_dma_dma_mem_ctl_dma_mem_write; // @[ifu.scala 129:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_wdata = io_ifu_dma_dma_mem_ctl_dma_mem_wdata; // @[ifu.scala 129:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_tag = io_ifu_dma_dma_mem_ctl_dma_mem_tag; // @[ifu.scala 129:26]
  assign mem_ctl_io_iccm_rd_data = io_iccm_rd_data; // @[ifu.scala 131:19]
  assign mem_ctl_io_iccm_rd_data_ecc = io_iccm_rd_data_ecc; // @[ifu.scala 131:19]
  assign mem_ctl_io_ic_rd_data = io_ic_rd_data; // @[ifu.scala 130:17]
  assign mem_ctl_io_ic_debug_rd_data = io_ic_debug_rd_data; // @[ifu.scala 130:17]
  assign mem_ctl_io_ic_tag_debug_rd_data = io_ic_tag_debug_rd_data; // @[ifu.scala 130:17]
  assign mem_ctl_io_ic_eccerr = io_ic_eccerr; // @[ifu.scala 130:17]
  assign mem_ctl_io_ic_rd_hit = io_ic_rd_hit; // @[ifu.scala 130:17]
  assign mem_ctl_io_ic_tag_perr = io_ic_tag_perr; // @[ifu.scala 130:17]
  assign mem_ctl_io_ifu_fetch_val = mem_ctl_io_ic_fetch_val_f; // @[ifu.scala 132:28]
  assign mem_ctl_io_dec_tlu_flush_lower_wb = io_dec_tlu_flush_lower_wb; // @[ifu.scala 133:37]
  assign bp_ctl_clock = clock;
  assign bp_ctl_reset = reset;
  assign bp_ctl_io_ic_hit_f = mem_ctl_io_ic_hit_f; // @[ifu.scala 104:22]
  assign bp_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 109:29]
  assign bp_ctl_io_ifc_fetch_addr_f = ifc_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 105:30]
  assign bp_ctl_io_ifc_fetch_req_f = ifc_ctl_io_ifc_fetch_req_f; // @[ifu.scala 106:29]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_valid = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid; // @[ifu.scala 107:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_hist = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist; // @[ifu.scala 107:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu.scala 107:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[ifu.scala 107:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_way = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu.scala 107:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_middle = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu.scala 107:20]
  assign bp_ctl_io_dec_bp_dec_tlu_flush_leak_one_wb = io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb; // @[ifu.scala 107:20]
  assign bp_ctl_io_dec_bp_dec_tlu_bpred_disable = io_ifu_dec_dec_bp_dec_tlu_bpred_disable; // @[ifu.scala 107:20]
  assign bp_ctl_io_dec_tlu_flush_lower_wb = io_dec_tlu_flush_lower_wb; // @[ifu.scala 110:36]
  assign bp_ctl_io_exu_bp_exu_i0_br_index_r = io_exu_ifu_exu_bp_exu_i0_br_index_r; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_i0_br_fghr_r = io_exu_ifu_exu_bp_exu_i0_br_fghr_r; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_valid = io_exu_ifu_exu_bp_exu_mp_pkt_valid; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_misp = io_exu_ifu_exu_bp_exu_mp_pkt_bits_misp; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_ataken = io_exu_ifu_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_boffset = io_exu_ifu_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pc4 = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pc4; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_hist = io_exu_ifu_exu_bp_exu_mp_pkt_bits_hist; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_toffset = io_exu_ifu_exu_bp_exu_mp_pkt_bits_toffset; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pcall = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pja = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pja; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_way = io_exu_ifu_exu_bp_exu_mp_pkt_bits_way; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pret = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pret; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_eghr = io_exu_ifu_exu_bp_exu_mp_eghr; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_fghr = io_exu_ifu_exu_bp_exu_mp_fghr; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_index = io_exu_ifu_exu_bp_exu_mp_index; // @[ifu.scala 108:20]
  assign bp_ctl_io_exu_bp_exu_mp_btag = io_exu_ifu_exu_bp_exu_mp_btag; // @[ifu.scala 108:20]
  assign aln_ctl_clk = clock;
  assign aln_ctl_reset = reset;
  assign aln_ctl_io_active_clk = io_active_clk; // @[ifu.scala 63:25]
  assign aln_ctl_io_ifu_async_error_start = mem_ctl_io_ifu_async_error_start; // @[ifu.scala 64:36]
  assign aln_ctl_io_iccm_rd_ecc_double_err = mem_ctl_io_iccm_rd_ecc_double_err; // @[ifu.scala 65:37]
  assign aln_ctl_io_ic_access_fault_f = mem_ctl_io_ic_access_fault_f; // @[ifu.scala 66:32]
  assign aln_ctl_io_ic_access_fault_type_f = mem_ctl_io_ic_access_fault_type_f; // @[ifu.scala 67:37]
  assign aln_ctl_io_dec_i0_decode_d = io_dec_i0_decode_d; // @[ifu.scala 94:30]
  assign aln_ctl_io_ifu_bp_fghr_f = bp_ctl_io_ifu_bp_fghr_f; // @[ifu.scala 68:28]
  assign aln_ctl_io_ifu_bp_btb_target_f = bp_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 69:34]
  assign aln_ctl_io_ifu_bp_poffset_f = bp_ctl_io_ifu_bp_poffset_f; // @[ifu.scala 70:31]
  assign aln_ctl_io_ifu_bp_hist0_f = bp_ctl_io_ifu_bp_hist0_f; // @[ifu.scala 71:29]
  assign aln_ctl_io_ifu_bp_hist1_f = bp_ctl_io_ifu_bp_hist1_f; // @[ifu.scala 72:29]
  assign aln_ctl_io_ifu_bp_pc4_f = bp_ctl_io_ifu_bp_pc4_f; // @[ifu.scala 73:27]
  assign aln_ctl_io_ifu_bp_way_f = bp_ctl_io_ifu_bp_way_f; // @[ifu.scala 74:27]
  assign aln_ctl_io_ifu_bp_valid_f = bp_ctl_io_ifu_bp_valid_f; // @[ifu.scala 75:29]
  assign aln_ctl_io_ifu_bp_ret_f = bp_ctl_io_ifu_bp_ret_f; // @[ifu.scala 76:27]
  assign aln_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 77:30]
  assign aln_ctl_io_ifu_fetch_data_f = mem_ctl_io_ic_data_f; // @[ifu.scala 97:31]
  assign aln_ctl_io_ifu_fetch_val = mem_ctl_io_ifu_fetch_val; // @[ifu.scala 98:28]
  assign aln_ctl_io_ifu_fetch_pc = ifc_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 99:27]
  assign ifc_ctl_clock = clock;
  assign ifc_ctl_reset = reset;
  assign ifc_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 52:30]
  assign ifc_ctl_io_exu_flush_path_final = io_exu_flush_path_final; // @[ifu.scala 59:35]
  assign ifc_ctl_io_free_l2clk = io_free_l2clk; // @[ifu.scala 46:25]
  assign ifc_ctl_io_ic_hit_f = mem_ctl_io_ic_hit_f; // @[ifu.scala 48:23]
  assign ifc_ctl_io_ifu_ic_mb_empty = mem_ctl_io_ifu_ic_mb_empty; // @[ifu.scala 58:30]
  assign ifc_ctl_io_ifu_fb_consume1 = aln_ctl_io_ifu_fb_consume1; // @[ifu.scala 49:30]
  assign ifc_ctl_io_ifu_fb_consume2 = aln_ctl_io_ifu_fb_consume2; // @[ifu.scala 50:30]
  assign ifc_ctl_io_ifu_bp_hit_taken_f = bp_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 53:33]
  assign ifc_ctl_io_ifu_bp_btb_target_f = bp_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 54:34]
  assign ifc_ctl_io_ic_dma_active = mem_ctl_io_ic_dma_active; // @[ifu.scala 55:28]
  assign ifc_ctl_io_ic_write_stall = mem_ctl_io_ic_write_stall; // @[ifu.scala 56:29]
  assign ifc_ctl_io_dec_ifc_dec_tlu_flush_noredir_wb = io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu.scala 51:22]
  assign ifc_ctl_io_dec_ifc_dec_tlu_mrac_ff = io_ifu_dec_dec_ifc_dec_tlu_mrac_ff; // @[ifu.scala 51:22]
  assign ifc_ctl_io_dma_ifc_dma_iccm_stall_any = io_ifu_dma_dma_ifc_dma_iccm_stall_any; // @[ifu.scala 57:22]
endmodule
