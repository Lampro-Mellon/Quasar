module el2_ifu_bp_ctl(
  input         clock,
  input         reset,
  input         io_active_clk,
  input         io_ic_hit_f,
  input  [30:0] io_ifc_fetch_addr_f,
  input         io_ifc_fetch_req_f,
  input         io_dec_tlu_br0_r_pkt_valid,
  input  [1:0]  io_dec_tlu_br0_r_pkt_hist,
  input         io_dec_tlu_br0_r_pkt_br_error,
  input         io_dec_tlu_br0_r_pkt_br_start_error,
  input         io_dec_tlu_br0_r_pkt_way,
  input         io_dec_tlu_br0_r_pkt_middle,
  input  [7:0]  io_exu_i0_br_fghr_r,
  input  [7:0]  io_exu_i0_br_index_r,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_leak_one_wb,
  input         io_dec_tlu_bpred_disable,
  input         io_exu_mp_pkt_misp,
  input         io_exu_mp_pkt_ataken,
  input         io_exu_mp_pkt_boffset,
  input         io_exu_mp_pkt_pc4,
  input  [1:0]  io_exu_mp_pkt_hist,
  input  [11:0] io_exu_mp_pkt_toffset,
  input         io_exu_mp_pkt_valid,
  input         io_exu_mp_pkt_br_error,
  input         io_exu_mp_pkt_br_start_error,
  input  [31:0] io_exu_mp_pkt_prett,
  input         io_exu_mp_pkt_pcall,
  input         io_exu_mp_pkt_pret,
  input         io_exu_mp_pkt_pja,
  input         io_exu_mp_pkt_way,
  input  [7:0]  io_exu_mp_eghr,
  input  [7:0]  io_exu_mp_fghr,
  input  [7:0]  io_exu_mp_index,
  input  [4:0]  io_exu_mp_btag,
  input         io_exu_flush_final,
  output        io_ifu_bp_hit_taken_f,
  output [30:0] io_ifu_bp_btb_target_f,
  output        io_ifu_bp_inst_mask_f,
  output [7:0]  io_ifu_bp_fghr_f,
  output [1:0]  io_ifu_bp_way_f,
  output [1:0]  io_ifu_bp_ret_f,
  output [1:0]  io_ifu_bp_hist1_f,
  output [1:0]  io_ifu_bp_hist0_f,
  output [1:0]  io_ifu_bp_pc4_f,
  output [1:0]  io_ifu_bp_valid_f,
  output [11:0] io_ifu_bp_poffset_f
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [255:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
`endif // RANDOMIZE_REG_INIT
  wire  _T_40 = io_dec_tlu_flush_leak_one_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_bp_ctl.scala 131:47]
  reg  leak_one_f_d1; // @[el2_ifu_bp_ctl.scala 125:56]
  wire  _T_41 = leak_one_f_d1 & io_dec_tlu_flush_lower_wb; // @[el2_ifu_bp_ctl.scala 131:93]
  wire  leak_one_f = _T_40 | _T_41; // @[el2_ifu_bp_ctl.scala 131:76]
  wire  _T = ~leak_one_f; // @[el2_ifu_bp_ctl.scala 70:46]
  wire  exu_mp_valid = io_exu_mp_pkt_misp & _T; // @[el2_ifu_bp_ctl.scala 70:44]
  wire  dec_tlu_error_wb = io_dec_tlu_br0_r_pkt_br_start_error | io_dec_tlu_br0_r_pkt_br_error; // @[el2_ifu_bp_ctl.scala 92:50]
  wire [7:0] _T_4 = io_ifc_fetch_addr_f[8:1] ^ io_ifc_fetch_addr_f[16:9]; // @[el2_lib.scala 186:46]
  wire [7:0] btb_rd_addr_f = _T_4 ^ io_ifc_fetch_addr_f[24:17]; // @[el2_lib.scala 186:84]
  wire [29:0] fetch_addr_p1_f = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[el2_ifu_bp_ctl.scala 100:51]
  wire [30:0] _T_8 = {fetch_addr_p1_f,1'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_11 = _T_8[8:1] ^ _T_8[16:9]; // @[el2_lib.scala 186:46]
  wire [7:0] btb_rd_addr_p1_f = _T_11 ^ _T_8[24:17]; // @[el2_lib.scala 186:84]
  wire  _T_143 = ~io_ifc_fetch_addr_f[0]; // @[el2_ifu_bp_ctl.scala 177:40]
  wire  _T_2108 = btb_rd_addr_f == 8'h0; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_0; // @[Reg.scala 27:20]
  wire [21:0] _T_2620 = _T_2108 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_2110 = btb_rd_addr_f == 8'h1; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_1; // @[Reg.scala 27:20]
  wire [21:0] _T_2621 = _T_2110 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2876 = _T_2620 | _T_2621; // @[Mux.scala 27:72]
  wire  _T_2112 = btb_rd_addr_f == 8'h2; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_2; // @[Reg.scala 27:20]
  wire [21:0] _T_2622 = _T_2112 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2877 = _T_2876 | _T_2622; // @[Mux.scala 27:72]
  wire  _T_2114 = btb_rd_addr_f == 8'h3; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_3; // @[Reg.scala 27:20]
  wire [21:0] _T_2623 = _T_2114 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2878 = _T_2877 | _T_2623; // @[Mux.scala 27:72]
  wire  _T_2116 = btb_rd_addr_f == 8'h4; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_4; // @[Reg.scala 27:20]
  wire [21:0] _T_2624 = _T_2116 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2879 = _T_2878 | _T_2624; // @[Mux.scala 27:72]
  wire  _T_2118 = btb_rd_addr_f == 8'h5; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_5; // @[Reg.scala 27:20]
  wire [21:0] _T_2625 = _T_2118 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2880 = _T_2879 | _T_2625; // @[Mux.scala 27:72]
  wire  _T_2120 = btb_rd_addr_f == 8'h6; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_6; // @[Reg.scala 27:20]
  wire [21:0] _T_2626 = _T_2120 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2881 = _T_2880 | _T_2626; // @[Mux.scala 27:72]
  wire  _T_2122 = btb_rd_addr_f == 8'h7; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_7; // @[Reg.scala 27:20]
  wire [21:0] _T_2627 = _T_2122 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2882 = _T_2881 | _T_2627; // @[Mux.scala 27:72]
  wire  _T_2124 = btb_rd_addr_f == 8'h8; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_8; // @[Reg.scala 27:20]
  wire [21:0] _T_2628 = _T_2124 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2883 = _T_2882 | _T_2628; // @[Mux.scala 27:72]
  wire  _T_2126 = btb_rd_addr_f == 8'h9; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_9; // @[Reg.scala 27:20]
  wire [21:0] _T_2629 = _T_2126 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2884 = _T_2883 | _T_2629; // @[Mux.scala 27:72]
  wire  _T_2128 = btb_rd_addr_f == 8'ha; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_10; // @[Reg.scala 27:20]
  wire [21:0] _T_2630 = _T_2128 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2885 = _T_2884 | _T_2630; // @[Mux.scala 27:72]
  wire  _T_2130 = btb_rd_addr_f == 8'hb; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_11; // @[Reg.scala 27:20]
  wire [21:0] _T_2631 = _T_2130 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2886 = _T_2885 | _T_2631; // @[Mux.scala 27:72]
  wire  _T_2132 = btb_rd_addr_f == 8'hc; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_12; // @[Reg.scala 27:20]
  wire [21:0] _T_2632 = _T_2132 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2887 = _T_2886 | _T_2632; // @[Mux.scala 27:72]
  wire  _T_2134 = btb_rd_addr_f == 8'hd; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_13; // @[Reg.scala 27:20]
  wire [21:0] _T_2633 = _T_2134 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2888 = _T_2887 | _T_2633; // @[Mux.scala 27:72]
  wire  _T_2136 = btb_rd_addr_f == 8'he; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_14; // @[Reg.scala 27:20]
  wire [21:0] _T_2634 = _T_2136 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2889 = _T_2888 | _T_2634; // @[Mux.scala 27:72]
  wire  _T_2138 = btb_rd_addr_f == 8'hf; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_15; // @[Reg.scala 27:20]
  wire [21:0] _T_2635 = _T_2138 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2890 = _T_2889 | _T_2635; // @[Mux.scala 27:72]
  wire  _T_2140 = btb_rd_addr_f == 8'h10; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_16; // @[Reg.scala 27:20]
  wire [21:0] _T_2636 = _T_2140 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2891 = _T_2890 | _T_2636; // @[Mux.scala 27:72]
  wire  _T_2142 = btb_rd_addr_f == 8'h11; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_17; // @[Reg.scala 27:20]
  wire [21:0] _T_2637 = _T_2142 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2892 = _T_2891 | _T_2637; // @[Mux.scala 27:72]
  wire  _T_2144 = btb_rd_addr_f == 8'h12; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_18; // @[Reg.scala 27:20]
  wire [21:0] _T_2638 = _T_2144 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2893 = _T_2892 | _T_2638; // @[Mux.scala 27:72]
  wire  _T_2146 = btb_rd_addr_f == 8'h13; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_19; // @[Reg.scala 27:20]
  wire [21:0] _T_2639 = _T_2146 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2894 = _T_2893 | _T_2639; // @[Mux.scala 27:72]
  wire  _T_2148 = btb_rd_addr_f == 8'h14; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_20; // @[Reg.scala 27:20]
  wire [21:0] _T_2640 = _T_2148 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2895 = _T_2894 | _T_2640; // @[Mux.scala 27:72]
  wire  _T_2150 = btb_rd_addr_f == 8'h15; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_21; // @[Reg.scala 27:20]
  wire [21:0] _T_2641 = _T_2150 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2896 = _T_2895 | _T_2641; // @[Mux.scala 27:72]
  wire  _T_2152 = btb_rd_addr_f == 8'h16; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_22; // @[Reg.scala 27:20]
  wire [21:0] _T_2642 = _T_2152 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2897 = _T_2896 | _T_2642; // @[Mux.scala 27:72]
  wire  _T_2154 = btb_rd_addr_f == 8'h17; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_23; // @[Reg.scala 27:20]
  wire [21:0] _T_2643 = _T_2154 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2898 = _T_2897 | _T_2643; // @[Mux.scala 27:72]
  wire  _T_2156 = btb_rd_addr_f == 8'h18; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_24; // @[Reg.scala 27:20]
  wire [21:0] _T_2644 = _T_2156 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2899 = _T_2898 | _T_2644; // @[Mux.scala 27:72]
  wire  _T_2158 = btb_rd_addr_f == 8'h19; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_25; // @[Reg.scala 27:20]
  wire [21:0] _T_2645 = _T_2158 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2900 = _T_2899 | _T_2645; // @[Mux.scala 27:72]
  wire  _T_2160 = btb_rd_addr_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_26; // @[Reg.scala 27:20]
  wire [21:0] _T_2646 = _T_2160 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2901 = _T_2900 | _T_2646; // @[Mux.scala 27:72]
  wire  _T_2162 = btb_rd_addr_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_27; // @[Reg.scala 27:20]
  wire [21:0] _T_2647 = _T_2162 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2902 = _T_2901 | _T_2647; // @[Mux.scala 27:72]
  wire  _T_2164 = btb_rd_addr_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_28; // @[Reg.scala 27:20]
  wire [21:0] _T_2648 = _T_2164 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2903 = _T_2902 | _T_2648; // @[Mux.scala 27:72]
  wire  _T_2166 = btb_rd_addr_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_29; // @[Reg.scala 27:20]
  wire [21:0] _T_2649 = _T_2166 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2904 = _T_2903 | _T_2649; // @[Mux.scala 27:72]
  wire  _T_2168 = btb_rd_addr_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_30; // @[Reg.scala 27:20]
  wire [21:0] _T_2650 = _T_2168 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2905 = _T_2904 | _T_2650; // @[Mux.scala 27:72]
  wire  _T_2170 = btb_rd_addr_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_31; // @[Reg.scala 27:20]
  wire [21:0] _T_2651 = _T_2170 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2906 = _T_2905 | _T_2651; // @[Mux.scala 27:72]
  wire  _T_2172 = btb_rd_addr_f == 8'h20; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_32; // @[Reg.scala 27:20]
  wire [21:0] _T_2652 = _T_2172 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2907 = _T_2906 | _T_2652; // @[Mux.scala 27:72]
  wire  _T_2174 = btb_rd_addr_f == 8'h21; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_33; // @[Reg.scala 27:20]
  wire [21:0] _T_2653 = _T_2174 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2908 = _T_2907 | _T_2653; // @[Mux.scala 27:72]
  wire  _T_2176 = btb_rd_addr_f == 8'h22; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_34; // @[Reg.scala 27:20]
  wire [21:0] _T_2654 = _T_2176 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2909 = _T_2908 | _T_2654; // @[Mux.scala 27:72]
  wire  _T_2178 = btb_rd_addr_f == 8'h23; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_35; // @[Reg.scala 27:20]
  wire [21:0] _T_2655 = _T_2178 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2910 = _T_2909 | _T_2655; // @[Mux.scala 27:72]
  wire  _T_2180 = btb_rd_addr_f == 8'h24; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_36; // @[Reg.scala 27:20]
  wire [21:0] _T_2656 = _T_2180 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2911 = _T_2910 | _T_2656; // @[Mux.scala 27:72]
  wire  _T_2182 = btb_rd_addr_f == 8'h25; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_37; // @[Reg.scala 27:20]
  wire [21:0] _T_2657 = _T_2182 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2912 = _T_2911 | _T_2657; // @[Mux.scala 27:72]
  wire  _T_2184 = btb_rd_addr_f == 8'h26; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_38; // @[Reg.scala 27:20]
  wire [21:0] _T_2658 = _T_2184 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2913 = _T_2912 | _T_2658; // @[Mux.scala 27:72]
  wire  _T_2186 = btb_rd_addr_f == 8'h27; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_39; // @[Reg.scala 27:20]
  wire [21:0] _T_2659 = _T_2186 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2914 = _T_2913 | _T_2659; // @[Mux.scala 27:72]
  wire  _T_2188 = btb_rd_addr_f == 8'h28; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_40; // @[Reg.scala 27:20]
  wire [21:0] _T_2660 = _T_2188 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2915 = _T_2914 | _T_2660; // @[Mux.scala 27:72]
  wire  _T_2190 = btb_rd_addr_f == 8'h29; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_41; // @[Reg.scala 27:20]
  wire [21:0] _T_2661 = _T_2190 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2916 = _T_2915 | _T_2661; // @[Mux.scala 27:72]
  wire  _T_2192 = btb_rd_addr_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_42; // @[Reg.scala 27:20]
  wire [21:0] _T_2662 = _T_2192 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2917 = _T_2916 | _T_2662; // @[Mux.scala 27:72]
  wire  _T_2194 = btb_rd_addr_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_43; // @[Reg.scala 27:20]
  wire [21:0] _T_2663 = _T_2194 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2918 = _T_2917 | _T_2663; // @[Mux.scala 27:72]
  wire  _T_2196 = btb_rd_addr_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_44; // @[Reg.scala 27:20]
  wire [21:0] _T_2664 = _T_2196 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2919 = _T_2918 | _T_2664; // @[Mux.scala 27:72]
  wire  _T_2198 = btb_rd_addr_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_45; // @[Reg.scala 27:20]
  wire [21:0] _T_2665 = _T_2198 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2920 = _T_2919 | _T_2665; // @[Mux.scala 27:72]
  wire  _T_2200 = btb_rd_addr_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_46; // @[Reg.scala 27:20]
  wire [21:0] _T_2666 = _T_2200 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2921 = _T_2920 | _T_2666; // @[Mux.scala 27:72]
  wire  _T_2202 = btb_rd_addr_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_47; // @[Reg.scala 27:20]
  wire [21:0] _T_2667 = _T_2202 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2922 = _T_2921 | _T_2667; // @[Mux.scala 27:72]
  wire  _T_2204 = btb_rd_addr_f == 8'h30; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_48; // @[Reg.scala 27:20]
  wire [21:0] _T_2668 = _T_2204 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2923 = _T_2922 | _T_2668; // @[Mux.scala 27:72]
  wire  _T_2206 = btb_rd_addr_f == 8'h31; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_49; // @[Reg.scala 27:20]
  wire [21:0] _T_2669 = _T_2206 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2924 = _T_2923 | _T_2669; // @[Mux.scala 27:72]
  wire  _T_2208 = btb_rd_addr_f == 8'h32; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_50; // @[Reg.scala 27:20]
  wire [21:0] _T_2670 = _T_2208 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2925 = _T_2924 | _T_2670; // @[Mux.scala 27:72]
  wire  _T_2210 = btb_rd_addr_f == 8'h33; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_51; // @[Reg.scala 27:20]
  wire [21:0] _T_2671 = _T_2210 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2926 = _T_2925 | _T_2671; // @[Mux.scala 27:72]
  wire  _T_2212 = btb_rd_addr_f == 8'h34; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_52; // @[Reg.scala 27:20]
  wire [21:0] _T_2672 = _T_2212 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2927 = _T_2926 | _T_2672; // @[Mux.scala 27:72]
  wire  _T_2214 = btb_rd_addr_f == 8'h35; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_53; // @[Reg.scala 27:20]
  wire [21:0] _T_2673 = _T_2214 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2928 = _T_2927 | _T_2673; // @[Mux.scala 27:72]
  wire  _T_2216 = btb_rd_addr_f == 8'h36; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_54; // @[Reg.scala 27:20]
  wire [21:0] _T_2674 = _T_2216 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2929 = _T_2928 | _T_2674; // @[Mux.scala 27:72]
  wire  _T_2218 = btb_rd_addr_f == 8'h37; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_55; // @[Reg.scala 27:20]
  wire [21:0] _T_2675 = _T_2218 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2930 = _T_2929 | _T_2675; // @[Mux.scala 27:72]
  wire  _T_2220 = btb_rd_addr_f == 8'h38; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_56; // @[Reg.scala 27:20]
  wire [21:0] _T_2676 = _T_2220 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2931 = _T_2930 | _T_2676; // @[Mux.scala 27:72]
  wire  _T_2222 = btb_rd_addr_f == 8'h39; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_57; // @[Reg.scala 27:20]
  wire [21:0] _T_2677 = _T_2222 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2932 = _T_2931 | _T_2677; // @[Mux.scala 27:72]
  wire  _T_2224 = btb_rd_addr_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_58; // @[Reg.scala 27:20]
  wire [21:0] _T_2678 = _T_2224 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2933 = _T_2932 | _T_2678; // @[Mux.scala 27:72]
  wire  _T_2226 = btb_rd_addr_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_59; // @[Reg.scala 27:20]
  wire [21:0] _T_2679 = _T_2226 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2934 = _T_2933 | _T_2679; // @[Mux.scala 27:72]
  wire  _T_2228 = btb_rd_addr_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_60; // @[Reg.scala 27:20]
  wire [21:0] _T_2680 = _T_2228 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2935 = _T_2934 | _T_2680; // @[Mux.scala 27:72]
  wire  _T_2230 = btb_rd_addr_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_61; // @[Reg.scala 27:20]
  wire [21:0] _T_2681 = _T_2230 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2936 = _T_2935 | _T_2681; // @[Mux.scala 27:72]
  wire  _T_2232 = btb_rd_addr_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_62; // @[Reg.scala 27:20]
  wire [21:0] _T_2682 = _T_2232 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2937 = _T_2936 | _T_2682; // @[Mux.scala 27:72]
  wire  _T_2234 = btb_rd_addr_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_63; // @[Reg.scala 27:20]
  wire [21:0] _T_2683 = _T_2234 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2938 = _T_2937 | _T_2683; // @[Mux.scala 27:72]
  wire  _T_2236 = btb_rd_addr_f == 8'h40; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_64; // @[Reg.scala 27:20]
  wire [21:0] _T_2684 = _T_2236 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2939 = _T_2938 | _T_2684; // @[Mux.scala 27:72]
  wire  _T_2238 = btb_rd_addr_f == 8'h41; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_65; // @[Reg.scala 27:20]
  wire [21:0] _T_2685 = _T_2238 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2940 = _T_2939 | _T_2685; // @[Mux.scala 27:72]
  wire  _T_2240 = btb_rd_addr_f == 8'h42; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_66; // @[Reg.scala 27:20]
  wire [21:0] _T_2686 = _T_2240 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2941 = _T_2940 | _T_2686; // @[Mux.scala 27:72]
  wire  _T_2242 = btb_rd_addr_f == 8'h43; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_67; // @[Reg.scala 27:20]
  wire [21:0] _T_2687 = _T_2242 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2942 = _T_2941 | _T_2687; // @[Mux.scala 27:72]
  wire  _T_2244 = btb_rd_addr_f == 8'h44; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_68; // @[Reg.scala 27:20]
  wire [21:0] _T_2688 = _T_2244 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2943 = _T_2942 | _T_2688; // @[Mux.scala 27:72]
  wire  _T_2246 = btb_rd_addr_f == 8'h45; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_69; // @[Reg.scala 27:20]
  wire [21:0] _T_2689 = _T_2246 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2944 = _T_2943 | _T_2689; // @[Mux.scala 27:72]
  wire  _T_2248 = btb_rd_addr_f == 8'h46; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_70; // @[Reg.scala 27:20]
  wire [21:0] _T_2690 = _T_2248 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2945 = _T_2944 | _T_2690; // @[Mux.scala 27:72]
  wire  _T_2250 = btb_rd_addr_f == 8'h47; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_71; // @[Reg.scala 27:20]
  wire [21:0] _T_2691 = _T_2250 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2946 = _T_2945 | _T_2691; // @[Mux.scala 27:72]
  wire  _T_2252 = btb_rd_addr_f == 8'h48; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_72; // @[Reg.scala 27:20]
  wire [21:0] _T_2692 = _T_2252 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2947 = _T_2946 | _T_2692; // @[Mux.scala 27:72]
  wire  _T_2254 = btb_rd_addr_f == 8'h49; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_73; // @[Reg.scala 27:20]
  wire [21:0] _T_2693 = _T_2254 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2948 = _T_2947 | _T_2693; // @[Mux.scala 27:72]
  wire  _T_2256 = btb_rd_addr_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_74; // @[Reg.scala 27:20]
  wire [21:0] _T_2694 = _T_2256 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2949 = _T_2948 | _T_2694; // @[Mux.scala 27:72]
  wire  _T_2258 = btb_rd_addr_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_75; // @[Reg.scala 27:20]
  wire [21:0] _T_2695 = _T_2258 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2950 = _T_2949 | _T_2695; // @[Mux.scala 27:72]
  wire  _T_2260 = btb_rd_addr_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_76; // @[Reg.scala 27:20]
  wire [21:0] _T_2696 = _T_2260 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2951 = _T_2950 | _T_2696; // @[Mux.scala 27:72]
  wire  _T_2262 = btb_rd_addr_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_77; // @[Reg.scala 27:20]
  wire [21:0] _T_2697 = _T_2262 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2952 = _T_2951 | _T_2697; // @[Mux.scala 27:72]
  wire  _T_2264 = btb_rd_addr_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_78; // @[Reg.scala 27:20]
  wire [21:0] _T_2698 = _T_2264 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2953 = _T_2952 | _T_2698; // @[Mux.scala 27:72]
  wire  _T_2266 = btb_rd_addr_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_79; // @[Reg.scala 27:20]
  wire [21:0] _T_2699 = _T_2266 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2954 = _T_2953 | _T_2699; // @[Mux.scala 27:72]
  wire  _T_2268 = btb_rd_addr_f == 8'h50; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_80; // @[Reg.scala 27:20]
  wire [21:0] _T_2700 = _T_2268 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2955 = _T_2954 | _T_2700; // @[Mux.scala 27:72]
  wire  _T_2270 = btb_rd_addr_f == 8'h51; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_81; // @[Reg.scala 27:20]
  wire [21:0] _T_2701 = _T_2270 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2956 = _T_2955 | _T_2701; // @[Mux.scala 27:72]
  wire  _T_2272 = btb_rd_addr_f == 8'h52; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_82; // @[Reg.scala 27:20]
  wire [21:0] _T_2702 = _T_2272 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2957 = _T_2956 | _T_2702; // @[Mux.scala 27:72]
  wire  _T_2274 = btb_rd_addr_f == 8'h53; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_83; // @[Reg.scala 27:20]
  wire [21:0] _T_2703 = _T_2274 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2958 = _T_2957 | _T_2703; // @[Mux.scala 27:72]
  wire  _T_2276 = btb_rd_addr_f == 8'h54; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_84; // @[Reg.scala 27:20]
  wire [21:0] _T_2704 = _T_2276 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2959 = _T_2958 | _T_2704; // @[Mux.scala 27:72]
  wire  _T_2278 = btb_rd_addr_f == 8'h55; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_85; // @[Reg.scala 27:20]
  wire [21:0] _T_2705 = _T_2278 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2960 = _T_2959 | _T_2705; // @[Mux.scala 27:72]
  wire  _T_2280 = btb_rd_addr_f == 8'h56; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_86; // @[Reg.scala 27:20]
  wire [21:0] _T_2706 = _T_2280 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2961 = _T_2960 | _T_2706; // @[Mux.scala 27:72]
  wire  _T_2282 = btb_rd_addr_f == 8'h57; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_87; // @[Reg.scala 27:20]
  wire [21:0] _T_2707 = _T_2282 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2962 = _T_2961 | _T_2707; // @[Mux.scala 27:72]
  wire  _T_2284 = btb_rd_addr_f == 8'h58; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_88; // @[Reg.scala 27:20]
  wire [21:0] _T_2708 = _T_2284 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2963 = _T_2962 | _T_2708; // @[Mux.scala 27:72]
  wire  _T_2286 = btb_rd_addr_f == 8'h59; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_89; // @[Reg.scala 27:20]
  wire [21:0] _T_2709 = _T_2286 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2964 = _T_2963 | _T_2709; // @[Mux.scala 27:72]
  wire  _T_2288 = btb_rd_addr_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_90; // @[Reg.scala 27:20]
  wire [21:0] _T_2710 = _T_2288 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2965 = _T_2964 | _T_2710; // @[Mux.scala 27:72]
  wire  _T_2290 = btb_rd_addr_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_91; // @[Reg.scala 27:20]
  wire [21:0] _T_2711 = _T_2290 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2966 = _T_2965 | _T_2711; // @[Mux.scala 27:72]
  wire  _T_2292 = btb_rd_addr_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_92; // @[Reg.scala 27:20]
  wire [21:0] _T_2712 = _T_2292 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2967 = _T_2966 | _T_2712; // @[Mux.scala 27:72]
  wire  _T_2294 = btb_rd_addr_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_93; // @[Reg.scala 27:20]
  wire [21:0] _T_2713 = _T_2294 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2968 = _T_2967 | _T_2713; // @[Mux.scala 27:72]
  wire  _T_2296 = btb_rd_addr_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_94; // @[Reg.scala 27:20]
  wire [21:0] _T_2714 = _T_2296 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2969 = _T_2968 | _T_2714; // @[Mux.scala 27:72]
  wire  _T_2298 = btb_rd_addr_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_95; // @[Reg.scala 27:20]
  wire [21:0] _T_2715 = _T_2298 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2970 = _T_2969 | _T_2715; // @[Mux.scala 27:72]
  wire  _T_2300 = btb_rd_addr_f == 8'h60; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_96; // @[Reg.scala 27:20]
  wire [21:0] _T_2716 = _T_2300 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2971 = _T_2970 | _T_2716; // @[Mux.scala 27:72]
  wire  _T_2302 = btb_rd_addr_f == 8'h61; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_97; // @[Reg.scala 27:20]
  wire [21:0] _T_2717 = _T_2302 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2972 = _T_2971 | _T_2717; // @[Mux.scala 27:72]
  wire  _T_2304 = btb_rd_addr_f == 8'h62; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_98; // @[Reg.scala 27:20]
  wire [21:0] _T_2718 = _T_2304 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2973 = _T_2972 | _T_2718; // @[Mux.scala 27:72]
  wire  _T_2306 = btb_rd_addr_f == 8'h63; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_99; // @[Reg.scala 27:20]
  wire [21:0] _T_2719 = _T_2306 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2974 = _T_2973 | _T_2719; // @[Mux.scala 27:72]
  wire  _T_2308 = btb_rd_addr_f == 8'h64; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_100; // @[Reg.scala 27:20]
  wire [21:0] _T_2720 = _T_2308 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2975 = _T_2974 | _T_2720; // @[Mux.scala 27:72]
  wire  _T_2310 = btb_rd_addr_f == 8'h65; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_101; // @[Reg.scala 27:20]
  wire [21:0] _T_2721 = _T_2310 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2976 = _T_2975 | _T_2721; // @[Mux.scala 27:72]
  wire  _T_2312 = btb_rd_addr_f == 8'h66; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_102; // @[Reg.scala 27:20]
  wire [21:0] _T_2722 = _T_2312 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2977 = _T_2976 | _T_2722; // @[Mux.scala 27:72]
  wire  _T_2314 = btb_rd_addr_f == 8'h67; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_103; // @[Reg.scala 27:20]
  wire [21:0] _T_2723 = _T_2314 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2978 = _T_2977 | _T_2723; // @[Mux.scala 27:72]
  wire  _T_2316 = btb_rd_addr_f == 8'h68; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_104; // @[Reg.scala 27:20]
  wire [21:0] _T_2724 = _T_2316 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2979 = _T_2978 | _T_2724; // @[Mux.scala 27:72]
  wire  _T_2318 = btb_rd_addr_f == 8'h69; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_105; // @[Reg.scala 27:20]
  wire [21:0] _T_2725 = _T_2318 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2980 = _T_2979 | _T_2725; // @[Mux.scala 27:72]
  wire  _T_2320 = btb_rd_addr_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_106; // @[Reg.scala 27:20]
  wire [21:0] _T_2726 = _T_2320 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2981 = _T_2980 | _T_2726; // @[Mux.scala 27:72]
  wire  _T_2322 = btb_rd_addr_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_107; // @[Reg.scala 27:20]
  wire [21:0] _T_2727 = _T_2322 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2982 = _T_2981 | _T_2727; // @[Mux.scala 27:72]
  wire  _T_2324 = btb_rd_addr_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_108; // @[Reg.scala 27:20]
  wire [21:0] _T_2728 = _T_2324 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2983 = _T_2982 | _T_2728; // @[Mux.scala 27:72]
  wire  _T_2326 = btb_rd_addr_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_109; // @[Reg.scala 27:20]
  wire [21:0] _T_2729 = _T_2326 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2984 = _T_2983 | _T_2729; // @[Mux.scala 27:72]
  wire  _T_2328 = btb_rd_addr_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_110; // @[Reg.scala 27:20]
  wire [21:0] _T_2730 = _T_2328 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2985 = _T_2984 | _T_2730; // @[Mux.scala 27:72]
  wire  _T_2330 = btb_rd_addr_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_111; // @[Reg.scala 27:20]
  wire [21:0] _T_2731 = _T_2330 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2986 = _T_2985 | _T_2731; // @[Mux.scala 27:72]
  wire  _T_2332 = btb_rd_addr_f == 8'h70; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_112; // @[Reg.scala 27:20]
  wire [21:0] _T_2732 = _T_2332 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2987 = _T_2986 | _T_2732; // @[Mux.scala 27:72]
  wire  _T_2334 = btb_rd_addr_f == 8'h71; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_113; // @[Reg.scala 27:20]
  wire [21:0] _T_2733 = _T_2334 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2988 = _T_2987 | _T_2733; // @[Mux.scala 27:72]
  wire  _T_2336 = btb_rd_addr_f == 8'h72; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_114; // @[Reg.scala 27:20]
  wire [21:0] _T_2734 = _T_2336 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2989 = _T_2988 | _T_2734; // @[Mux.scala 27:72]
  wire  _T_2338 = btb_rd_addr_f == 8'h73; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_115; // @[Reg.scala 27:20]
  wire [21:0] _T_2735 = _T_2338 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2990 = _T_2989 | _T_2735; // @[Mux.scala 27:72]
  wire  _T_2340 = btb_rd_addr_f == 8'h74; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_116; // @[Reg.scala 27:20]
  wire [21:0] _T_2736 = _T_2340 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2991 = _T_2990 | _T_2736; // @[Mux.scala 27:72]
  wire  _T_2342 = btb_rd_addr_f == 8'h75; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_117; // @[Reg.scala 27:20]
  wire [21:0] _T_2737 = _T_2342 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2992 = _T_2991 | _T_2737; // @[Mux.scala 27:72]
  wire  _T_2344 = btb_rd_addr_f == 8'h76; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_118; // @[Reg.scala 27:20]
  wire [21:0] _T_2738 = _T_2344 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2993 = _T_2992 | _T_2738; // @[Mux.scala 27:72]
  wire  _T_2346 = btb_rd_addr_f == 8'h77; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_119; // @[Reg.scala 27:20]
  wire [21:0] _T_2739 = _T_2346 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2994 = _T_2993 | _T_2739; // @[Mux.scala 27:72]
  wire  _T_2348 = btb_rd_addr_f == 8'h78; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_120; // @[Reg.scala 27:20]
  wire [21:0] _T_2740 = _T_2348 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2995 = _T_2994 | _T_2740; // @[Mux.scala 27:72]
  wire  _T_2350 = btb_rd_addr_f == 8'h79; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_121; // @[Reg.scala 27:20]
  wire [21:0] _T_2741 = _T_2350 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2996 = _T_2995 | _T_2741; // @[Mux.scala 27:72]
  wire  _T_2352 = btb_rd_addr_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_122; // @[Reg.scala 27:20]
  wire [21:0] _T_2742 = _T_2352 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2997 = _T_2996 | _T_2742; // @[Mux.scala 27:72]
  wire  _T_2354 = btb_rd_addr_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_123; // @[Reg.scala 27:20]
  wire [21:0] _T_2743 = _T_2354 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2998 = _T_2997 | _T_2743; // @[Mux.scala 27:72]
  wire  _T_2356 = btb_rd_addr_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_124; // @[Reg.scala 27:20]
  wire [21:0] _T_2744 = _T_2356 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2999 = _T_2998 | _T_2744; // @[Mux.scala 27:72]
  wire  _T_2358 = btb_rd_addr_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_125; // @[Reg.scala 27:20]
  wire [21:0] _T_2745 = _T_2358 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3000 = _T_2999 | _T_2745; // @[Mux.scala 27:72]
  wire  _T_2360 = btb_rd_addr_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_126; // @[Reg.scala 27:20]
  wire [21:0] _T_2746 = _T_2360 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3001 = _T_3000 | _T_2746; // @[Mux.scala 27:72]
  wire  _T_2362 = btb_rd_addr_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_127; // @[Reg.scala 27:20]
  wire [21:0] _T_2747 = _T_2362 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3002 = _T_3001 | _T_2747; // @[Mux.scala 27:72]
  wire  _T_2364 = btb_rd_addr_f == 8'h80; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_128; // @[Reg.scala 27:20]
  wire [21:0] _T_2748 = _T_2364 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3003 = _T_3002 | _T_2748; // @[Mux.scala 27:72]
  wire  _T_2366 = btb_rd_addr_f == 8'h81; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_129; // @[Reg.scala 27:20]
  wire [21:0] _T_2749 = _T_2366 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3004 = _T_3003 | _T_2749; // @[Mux.scala 27:72]
  wire  _T_2368 = btb_rd_addr_f == 8'h82; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_130; // @[Reg.scala 27:20]
  wire [21:0] _T_2750 = _T_2368 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3005 = _T_3004 | _T_2750; // @[Mux.scala 27:72]
  wire  _T_2370 = btb_rd_addr_f == 8'h83; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_131; // @[Reg.scala 27:20]
  wire [21:0] _T_2751 = _T_2370 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3006 = _T_3005 | _T_2751; // @[Mux.scala 27:72]
  wire  _T_2372 = btb_rd_addr_f == 8'h84; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_132; // @[Reg.scala 27:20]
  wire [21:0] _T_2752 = _T_2372 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3007 = _T_3006 | _T_2752; // @[Mux.scala 27:72]
  wire  _T_2374 = btb_rd_addr_f == 8'h85; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_133; // @[Reg.scala 27:20]
  wire [21:0] _T_2753 = _T_2374 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3008 = _T_3007 | _T_2753; // @[Mux.scala 27:72]
  wire  _T_2376 = btb_rd_addr_f == 8'h86; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_134; // @[Reg.scala 27:20]
  wire [21:0] _T_2754 = _T_2376 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3009 = _T_3008 | _T_2754; // @[Mux.scala 27:72]
  wire  _T_2378 = btb_rd_addr_f == 8'h87; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_135; // @[Reg.scala 27:20]
  wire [21:0] _T_2755 = _T_2378 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3010 = _T_3009 | _T_2755; // @[Mux.scala 27:72]
  wire  _T_2380 = btb_rd_addr_f == 8'h88; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_136; // @[Reg.scala 27:20]
  wire [21:0] _T_2756 = _T_2380 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3011 = _T_3010 | _T_2756; // @[Mux.scala 27:72]
  wire  _T_2382 = btb_rd_addr_f == 8'h89; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_137; // @[Reg.scala 27:20]
  wire [21:0] _T_2757 = _T_2382 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3012 = _T_3011 | _T_2757; // @[Mux.scala 27:72]
  wire  _T_2384 = btb_rd_addr_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_138; // @[Reg.scala 27:20]
  wire [21:0] _T_2758 = _T_2384 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3013 = _T_3012 | _T_2758; // @[Mux.scala 27:72]
  wire  _T_2386 = btb_rd_addr_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_139; // @[Reg.scala 27:20]
  wire [21:0] _T_2759 = _T_2386 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3014 = _T_3013 | _T_2759; // @[Mux.scala 27:72]
  wire  _T_2388 = btb_rd_addr_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_140; // @[Reg.scala 27:20]
  wire [21:0] _T_2760 = _T_2388 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3015 = _T_3014 | _T_2760; // @[Mux.scala 27:72]
  wire  _T_2390 = btb_rd_addr_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_141; // @[Reg.scala 27:20]
  wire [21:0] _T_2761 = _T_2390 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3016 = _T_3015 | _T_2761; // @[Mux.scala 27:72]
  wire  _T_2392 = btb_rd_addr_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_142; // @[Reg.scala 27:20]
  wire [21:0] _T_2762 = _T_2392 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3017 = _T_3016 | _T_2762; // @[Mux.scala 27:72]
  wire  _T_2394 = btb_rd_addr_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_143; // @[Reg.scala 27:20]
  wire [21:0] _T_2763 = _T_2394 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3018 = _T_3017 | _T_2763; // @[Mux.scala 27:72]
  wire  _T_2396 = btb_rd_addr_f == 8'h90; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_144; // @[Reg.scala 27:20]
  wire [21:0] _T_2764 = _T_2396 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3019 = _T_3018 | _T_2764; // @[Mux.scala 27:72]
  wire  _T_2398 = btb_rd_addr_f == 8'h91; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_145; // @[Reg.scala 27:20]
  wire [21:0] _T_2765 = _T_2398 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3020 = _T_3019 | _T_2765; // @[Mux.scala 27:72]
  wire  _T_2400 = btb_rd_addr_f == 8'h92; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_146; // @[Reg.scala 27:20]
  wire [21:0] _T_2766 = _T_2400 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3021 = _T_3020 | _T_2766; // @[Mux.scala 27:72]
  wire  _T_2402 = btb_rd_addr_f == 8'h93; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_147; // @[Reg.scala 27:20]
  wire [21:0] _T_2767 = _T_2402 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3022 = _T_3021 | _T_2767; // @[Mux.scala 27:72]
  wire  _T_2404 = btb_rd_addr_f == 8'h94; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_148; // @[Reg.scala 27:20]
  wire [21:0] _T_2768 = _T_2404 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3023 = _T_3022 | _T_2768; // @[Mux.scala 27:72]
  wire  _T_2406 = btb_rd_addr_f == 8'h95; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_149; // @[Reg.scala 27:20]
  wire [21:0] _T_2769 = _T_2406 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3024 = _T_3023 | _T_2769; // @[Mux.scala 27:72]
  wire  _T_2408 = btb_rd_addr_f == 8'h96; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_150; // @[Reg.scala 27:20]
  wire [21:0] _T_2770 = _T_2408 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3025 = _T_3024 | _T_2770; // @[Mux.scala 27:72]
  wire  _T_2410 = btb_rd_addr_f == 8'h97; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_151; // @[Reg.scala 27:20]
  wire [21:0] _T_2771 = _T_2410 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3026 = _T_3025 | _T_2771; // @[Mux.scala 27:72]
  wire  _T_2412 = btb_rd_addr_f == 8'h98; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_152; // @[Reg.scala 27:20]
  wire [21:0] _T_2772 = _T_2412 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3027 = _T_3026 | _T_2772; // @[Mux.scala 27:72]
  wire  _T_2414 = btb_rd_addr_f == 8'h99; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_153; // @[Reg.scala 27:20]
  wire [21:0] _T_2773 = _T_2414 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3028 = _T_3027 | _T_2773; // @[Mux.scala 27:72]
  wire  _T_2416 = btb_rd_addr_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_154; // @[Reg.scala 27:20]
  wire [21:0] _T_2774 = _T_2416 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3029 = _T_3028 | _T_2774; // @[Mux.scala 27:72]
  wire  _T_2418 = btb_rd_addr_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_155; // @[Reg.scala 27:20]
  wire [21:0] _T_2775 = _T_2418 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3030 = _T_3029 | _T_2775; // @[Mux.scala 27:72]
  wire  _T_2420 = btb_rd_addr_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_156; // @[Reg.scala 27:20]
  wire [21:0] _T_2776 = _T_2420 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3031 = _T_3030 | _T_2776; // @[Mux.scala 27:72]
  wire  _T_2422 = btb_rd_addr_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_157; // @[Reg.scala 27:20]
  wire [21:0] _T_2777 = _T_2422 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3032 = _T_3031 | _T_2777; // @[Mux.scala 27:72]
  wire  _T_2424 = btb_rd_addr_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_158; // @[Reg.scala 27:20]
  wire [21:0] _T_2778 = _T_2424 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3033 = _T_3032 | _T_2778; // @[Mux.scala 27:72]
  wire  _T_2426 = btb_rd_addr_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_159; // @[Reg.scala 27:20]
  wire [21:0] _T_2779 = _T_2426 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3034 = _T_3033 | _T_2779; // @[Mux.scala 27:72]
  wire  _T_2428 = btb_rd_addr_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_160; // @[Reg.scala 27:20]
  wire [21:0] _T_2780 = _T_2428 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3035 = _T_3034 | _T_2780; // @[Mux.scala 27:72]
  wire  _T_2430 = btb_rd_addr_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_161; // @[Reg.scala 27:20]
  wire [21:0] _T_2781 = _T_2430 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3036 = _T_3035 | _T_2781; // @[Mux.scala 27:72]
  wire  _T_2432 = btb_rd_addr_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_162; // @[Reg.scala 27:20]
  wire [21:0] _T_2782 = _T_2432 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3037 = _T_3036 | _T_2782; // @[Mux.scala 27:72]
  wire  _T_2434 = btb_rd_addr_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_163; // @[Reg.scala 27:20]
  wire [21:0] _T_2783 = _T_2434 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3038 = _T_3037 | _T_2783; // @[Mux.scala 27:72]
  wire  _T_2436 = btb_rd_addr_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_164; // @[Reg.scala 27:20]
  wire [21:0] _T_2784 = _T_2436 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3039 = _T_3038 | _T_2784; // @[Mux.scala 27:72]
  wire  _T_2438 = btb_rd_addr_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_165; // @[Reg.scala 27:20]
  wire [21:0] _T_2785 = _T_2438 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3040 = _T_3039 | _T_2785; // @[Mux.scala 27:72]
  wire  _T_2440 = btb_rd_addr_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_166; // @[Reg.scala 27:20]
  wire [21:0] _T_2786 = _T_2440 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3041 = _T_3040 | _T_2786; // @[Mux.scala 27:72]
  wire  _T_2442 = btb_rd_addr_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_167; // @[Reg.scala 27:20]
  wire [21:0] _T_2787 = _T_2442 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3042 = _T_3041 | _T_2787; // @[Mux.scala 27:72]
  wire  _T_2444 = btb_rd_addr_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_168; // @[Reg.scala 27:20]
  wire [21:0] _T_2788 = _T_2444 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3043 = _T_3042 | _T_2788; // @[Mux.scala 27:72]
  wire  _T_2446 = btb_rd_addr_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_169; // @[Reg.scala 27:20]
  wire [21:0] _T_2789 = _T_2446 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3044 = _T_3043 | _T_2789; // @[Mux.scala 27:72]
  wire  _T_2448 = btb_rd_addr_f == 8'haa; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_170; // @[Reg.scala 27:20]
  wire [21:0] _T_2790 = _T_2448 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3045 = _T_3044 | _T_2790; // @[Mux.scala 27:72]
  wire  _T_2450 = btb_rd_addr_f == 8'hab; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_171; // @[Reg.scala 27:20]
  wire [21:0] _T_2791 = _T_2450 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3046 = _T_3045 | _T_2791; // @[Mux.scala 27:72]
  wire  _T_2452 = btb_rd_addr_f == 8'hac; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_172; // @[Reg.scala 27:20]
  wire [21:0] _T_2792 = _T_2452 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3047 = _T_3046 | _T_2792; // @[Mux.scala 27:72]
  wire  _T_2454 = btb_rd_addr_f == 8'had; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_173; // @[Reg.scala 27:20]
  wire [21:0] _T_2793 = _T_2454 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3048 = _T_3047 | _T_2793; // @[Mux.scala 27:72]
  wire  _T_2456 = btb_rd_addr_f == 8'hae; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_174; // @[Reg.scala 27:20]
  wire [21:0] _T_2794 = _T_2456 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3049 = _T_3048 | _T_2794; // @[Mux.scala 27:72]
  wire  _T_2458 = btb_rd_addr_f == 8'haf; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_175; // @[Reg.scala 27:20]
  wire [21:0] _T_2795 = _T_2458 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3050 = _T_3049 | _T_2795; // @[Mux.scala 27:72]
  wire  _T_2460 = btb_rd_addr_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_176; // @[Reg.scala 27:20]
  wire [21:0] _T_2796 = _T_2460 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3051 = _T_3050 | _T_2796; // @[Mux.scala 27:72]
  wire  _T_2462 = btb_rd_addr_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_177; // @[Reg.scala 27:20]
  wire [21:0] _T_2797 = _T_2462 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3052 = _T_3051 | _T_2797; // @[Mux.scala 27:72]
  wire  _T_2464 = btb_rd_addr_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_178; // @[Reg.scala 27:20]
  wire [21:0] _T_2798 = _T_2464 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3053 = _T_3052 | _T_2798; // @[Mux.scala 27:72]
  wire  _T_2466 = btb_rd_addr_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_179; // @[Reg.scala 27:20]
  wire [21:0] _T_2799 = _T_2466 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3054 = _T_3053 | _T_2799; // @[Mux.scala 27:72]
  wire  _T_2468 = btb_rd_addr_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_180; // @[Reg.scala 27:20]
  wire [21:0] _T_2800 = _T_2468 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3055 = _T_3054 | _T_2800; // @[Mux.scala 27:72]
  wire  _T_2470 = btb_rd_addr_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_181; // @[Reg.scala 27:20]
  wire [21:0] _T_2801 = _T_2470 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3056 = _T_3055 | _T_2801; // @[Mux.scala 27:72]
  wire  _T_2472 = btb_rd_addr_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_182; // @[Reg.scala 27:20]
  wire [21:0] _T_2802 = _T_2472 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3057 = _T_3056 | _T_2802; // @[Mux.scala 27:72]
  wire  _T_2474 = btb_rd_addr_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_183; // @[Reg.scala 27:20]
  wire [21:0] _T_2803 = _T_2474 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3058 = _T_3057 | _T_2803; // @[Mux.scala 27:72]
  wire  _T_2476 = btb_rd_addr_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_184; // @[Reg.scala 27:20]
  wire [21:0] _T_2804 = _T_2476 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3059 = _T_3058 | _T_2804; // @[Mux.scala 27:72]
  wire  _T_2478 = btb_rd_addr_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_185; // @[Reg.scala 27:20]
  wire [21:0] _T_2805 = _T_2478 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3060 = _T_3059 | _T_2805; // @[Mux.scala 27:72]
  wire  _T_2480 = btb_rd_addr_f == 8'hba; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_186; // @[Reg.scala 27:20]
  wire [21:0] _T_2806 = _T_2480 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3061 = _T_3060 | _T_2806; // @[Mux.scala 27:72]
  wire  _T_2482 = btb_rd_addr_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_187; // @[Reg.scala 27:20]
  wire [21:0] _T_2807 = _T_2482 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3062 = _T_3061 | _T_2807; // @[Mux.scala 27:72]
  wire  _T_2484 = btb_rd_addr_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_188; // @[Reg.scala 27:20]
  wire [21:0] _T_2808 = _T_2484 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3063 = _T_3062 | _T_2808; // @[Mux.scala 27:72]
  wire  _T_2486 = btb_rd_addr_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_189; // @[Reg.scala 27:20]
  wire [21:0] _T_2809 = _T_2486 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3064 = _T_3063 | _T_2809; // @[Mux.scala 27:72]
  wire  _T_2488 = btb_rd_addr_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_190; // @[Reg.scala 27:20]
  wire [21:0] _T_2810 = _T_2488 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3065 = _T_3064 | _T_2810; // @[Mux.scala 27:72]
  wire  _T_2490 = btb_rd_addr_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_191; // @[Reg.scala 27:20]
  wire [21:0] _T_2811 = _T_2490 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3066 = _T_3065 | _T_2811; // @[Mux.scala 27:72]
  wire  _T_2492 = btb_rd_addr_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_192; // @[Reg.scala 27:20]
  wire [21:0] _T_2812 = _T_2492 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3067 = _T_3066 | _T_2812; // @[Mux.scala 27:72]
  wire  _T_2494 = btb_rd_addr_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_193; // @[Reg.scala 27:20]
  wire [21:0] _T_2813 = _T_2494 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3068 = _T_3067 | _T_2813; // @[Mux.scala 27:72]
  wire  _T_2496 = btb_rd_addr_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_194; // @[Reg.scala 27:20]
  wire [21:0] _T_2814 = _T_2496 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3069 = _T_3068 | _T_2814; // @[Mux.scala 27:72]
  wire  _T_2498 = btb_rd_addr_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_195; // @[Reg.scala 27:20]
  wire [21:0] _T_2815 = _T_2498 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3070 = _T_3069 | _T_2815; // @[Mux.scala 27:72]
  wire  _T_2500 = btb_rd_addr_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_196; // @[Reg.scala 27:20]
  wire [21:0] _T_2816 = _T_2500 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3071 = _T_3070 | _T_2816; // @[Mux.scala 27:72]
  wire  _T_2502 = btb_rd_addr_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_197; // @[Reg.scala 27:20]
  wire [21:0] _T_2817 = _T_2502 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3072 = _T_3071 | _T_2817; // @[Mux.scala 27:72]
  wire  _T_2504 = btb_rd_addr_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_198; // @[Reg.scala 27:20]
  wire [21:0] _T_2818 = _T_2504 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3073 = _T_3072 | _T_2818; // @[Mux.scala 27:72]
  wire  _T_2506 = btb_rd_addr_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_199; // @[Reg.scala 27:20]
  wire [21:0] _T_2819 = _T_2506 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3074 = _T_3073 | _T_2819; // @[Mux.scala 27:72]
  wire  _T_2508 = btb_rd_addr_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_200; // @[Reg.scala 27:20]
  wire [21:0] _T_2820 = _T_2508 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3075 = _T_3074 | _T_2820; // @[Mux.scala 27:72]
  wire  _T_2510 = btb_rd_addr_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_201; // @[Reg.scala 27:20]
  wire [21:0] _T_2821 = _T_2510 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3076 = _T_3075 | _T_2821; // @[Mux.scala 27:72]
  wire  _T_2512 = btb_rd_addr_f == 8'hca; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_202; // @[Reg.scala 27:20]
  wire [21:0] _T_2822 = _T_2512 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3077 = _T_3076 | _T_2822; // @[Mux.scala 27:72]
  wire  _T_2514 = btb_rd_addr_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_203; // @[Reg.scala 27:20]
  wire [21:0] _T_2823 = _T_2514 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3078 = _T_3077 | _T_2823; // @[Mux.scala 27:72]
  wire  _T_2516 = btb_rd_addr_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_204; // @[Reg.scala 27:20]
  wire [21:0] _T_2824 = _T_2516 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3079 = _T_3078 | _T_2824; // @[Mux.scala 27:72]
  wire  _T_2518 = btb_rd_addr_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_205; // @[Reg.scala 27:20]
  wire [21:0] _T_2825 = _T_2518 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3080 = _T_3079 | _T_2825; // @[Mux.scala 27:72]
  wire  _T_2520 = btb_rd_addr_f == 8'hce; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_206; // @[Reg.scala 27:20]
  wire [21:0] _T_2826 = _T_2520 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3081 = _T_3080 | _T_2826; // @[Mux.scala 27:72]
  wire  _T_2522 = btb_rd_addr_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_207; // @[Reg.scala 27:20]
  wire [21:0] _T_2827 = _T_2522 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3082 = _T_3081 | _T_2827; // @[Mux.scala 27:72]
  wire  _T_2524 = btb_rd_addr_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_208; // @[Reg.scala 27:20]
  wire [21:0] _T_2828 = _T_2524 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3083 = _T_3082 | _T_2828; // @[Mux.scala 27:72]
  wire  _T_2526 = btb_rd_addr_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_209; // @[Reg.scala 27:20]
  wire [21:0] _T_2829 = _T_2526 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3084 = _T_3083 | _T_2829; // @[Mux.scala 27:72]
  wire  _T_2528 = btb_rd_addr_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_210; // @[Reg.scala 27:20]
  wire [21:0] _T_2830 = _T_2528 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3085 = _T_3084 | _T_2830; // @[Mux.scala 27:72]
  wire  _T_2530 = btb_rd_addr_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_211; // @[Reg.scala 27:20]
  wire [21:0] _T_2831 = _T_2530 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3086 = _T_3085 | _T_2831; // @[Mux.scala 27:72]
  wire  _T_2532 = btb_rd_addr_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_212; // @[Reg.scala 27:20]
  wire [21:0] _T_2832 = _T_2532 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3087 = _T_3086 | _T_2832; // @[Mux.scala 27:72]
  wire  _T_2534 = btb_rd_addr_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_213; // @[Reg.scala 27:20]
  wire [21:0] _T_2833 = _T_2534 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3088 = _T_3087 | _T_2833; // @[Mux.scala 27:72]
  wire  _T_2536 = btb_rd_addr_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_214; // @[Reg.scala 27:20]
  wire [21:0] _T_2834 = _T_2536 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3089 = _T_3088 | _T_2834; // @[Mux.scala 27:72]
  wire  _T_2538 = btb_rd_addr_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_215; // @[Reg.scala 27:20]
  wire [21:0] _T_2835 = _T_2538 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3090 = _T_3089 | _T_2835; // @[Mux.scala 27:72]
  wire  _T_2540 = btb_rd_addr_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_216; // @[Reg.scala 27:20]
  wire [21:0] _T_2836 = _T_2540 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3091 = _T_3090 | _T_2836; // @[Mux.scala 27:72]
  wire  _T_2542 = btb_rd_addr_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_217; // @[Reg.scala 27:20]
  wire [21:0] _T_2837 = _T_2542 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3092 = _T_3091 | _T_2837; // @[Mux.scala 27:72]
  wire  _T_2544 = btb_rd_addr_f == 8'hda; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_218; // @[Reg.scala 27:20]
  wire [21:0] _T_2838 = _T_2544 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3093 = _T_3092 | _T_2838; // @[Mux.scala 27:72]
  wire  _T_2546 = btb_rd_addr_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_219; // @[Reg.scala 27:20]
  wire [21:0] _T_2839 = _T_2546 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3094 = _T_3093 | _T_2839; // @[Mux.scala 27:72]
  wire  _T_2548 = btb_rd_addr_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_220; // @[Reg.scala 27:20]
  wire [21:0] _T_2840 = _T_2548 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3095 = _T_3094 | _T_2840; // @[Mux.scala 27:72]
  wire  _T_2550 = btb_rd_addr_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_221; // @[Reg.scala 27:20]
  wire [21:0] _T_2841 = _T_2550 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3096 = _T_3095 | _T_2841; // @[Mux.scala 27:72]
  wire  _T_2552 = btb_rd_addr_f == 8'hde; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_222; // @[Reg.scala 27:20]
  wire [21:0] _T_2842 = _T_2552 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3097 = _T_3096 | _T_2842; // @[Mux.scala 27:72]
  wire  _T_2554 = btb_rd_addr_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_223; // @[Reg.scala 27:20]
  wire [21:0] _T_2843 = _T_2554 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3098 = _T_3097 | _T_2843; // @[Mux.scala 27:72]
  wire  _T_2556 = btb_rd_addr_f == 8'he0; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_224; // @[Reg.scala 27:20]
  wire [21:0] _T_2844 = _T_2556 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3099 = _T_3098 | _T_2844; // @[Mux.scala 27:72]
  wire  _T_2558 = btb_rd_addr_f == 8'he1; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_225; // @[Reg.scala 27:20]
  wire [21:0] _T_2845 = _T_2558 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3100 = _T_3099 | _T_2845; // @[Mux.scala 27:72]
  wire  _T_2560 = btb_rd_addr_f == 8'he2; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_226; // @[Reg.scala 27:20]
  wire [21:0] _T_2846 = _T_2560 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3101 = _T_3100 | _T_2846; // @[Mux.scala 27:72]
  wire  _T_2562 = btb_rd_addr_f == 8'he3; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_227; // @[Reg.scala 27:20]
  wire [21:0] _T_2847 = _T_2562 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3102 = _T_3101 | _T_2847; // @[Mux.scala 27:72]
  wire  _T_2564 = btb_rd_addr_f == 8'he4; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_228; // @[Reg.scala 27:20]
  wire [21:0] _T_2848 = _T_2564 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3103 = _T_3102 | _T_2848; // @[Mux.scala 27:72]
  wire  _T_2566 = btb_rd_addr_f == 8'he5; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_229; // @[Reg.scala 27:20]
  wire [21:0] _T_2849 = _T_2566 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3104 = _T_3103 | _T_2849; // @[Mux.scala 27:72]
  wire  _T_2568 = btb_rd_addr_f == 8'he6; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_230; // @[Reg.scala 27:20]
  wire [21:0] _T_2850 = _T_2568 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3105 = _T_3104 | _T_2850; // @[Mux.scala 27:72]
  wire  _T_2570 = btb_rd_addr_f == 8'he7; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_231; // @[Reg.scala 27:20]
  wire [21:0] _T_2851 = _T_2570 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3106 = _T_3105 | _T_2851; // @[Mux.scala 27:72]
  wire  _T_2572 = btb_rd_addr_f == 8'he8; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_232; // @[Reg.scala 27:20]
  wire [21:0] _T_2852 = _T_2572 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3107 = _T_3106 | _T_2852; // @[Mux.scala 27:72]
  wire  _T_2574 = btb_rd_addr_f == 8'he9; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_233; // @[Reg.scala 27:20]
  wire [21:0] _T_2853 = _T_2574 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3108 = _T_3107 | _T_2853; // @[Mux.scala 27:72]
  wire  _T_2576 = btb_rd_addr_f == 8'hea; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_234; // @[Reg.scala 27:20]
  wire [21:0] _T_2854 = _T_2576 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3109 = _T_3108 | _T_2854; // @[Mux.scala 27:72]
  wire  _T_2578 = btb_rd_addr_f == 8'heb; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_235; // @[Reg.scala 27:20]
  wire [21:0] _T_2855 = _T_2578 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3110 = _T_3109 | _T_2855; // @[Mux.scala 27:72]
  wire  _T_2580 = btb_rd_addr_f == 8'hec; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_236; // @[Reg.scala 27:20]
  wire [21:0] _T_2856 = _T_2580 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3111 = _T_3110 | _T_2856; // @[Mux.scala 27:72]
  wire  _T_2582 = btb_rd_addr_f == 8'hed; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_237; // @[Reg.scala 27:20]
  wire [21:0] _T_2857 = _T_2582 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3112 = _T_3111 | _T_2857; // @[Mux.scala 27:72]
  wire  _T_2584 = btb_rd_addr_f == 8'hee; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_238; // @[Reg.scala 27:20]
  wire [21:0] _T_2858 = _T_2584 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3113 = _T_3112 | _T_2858; // @[Mux.scala 27:72]
  wire  _T_2586 = btb_rd_addr_f == 8'hef; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_239; // @[Reg.scala 27:20]
  wire [21:0] _T_2859 = _T_2586 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3114 = _T_3113 | _T_2859; // @[Mux.scala 27:72]
  wire  _T_2588 = btb_rd_addr_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_240; // @[Reg.scala 27:20]
  wire [21:0] _T_2860 = _T_2588 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3115 = _T_3114 | _T_2860; // @[Mux.scala 27:72]
  wire  _T_2590 = btb_rd_addr_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_241; // @[Reg.scala 27:20]
  wire [21:0] _T_2861 = _T_2590 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3116 = _T_3115 | _T_2861; // @[Mux.scala 27:72]
  wire  _T_2592 = btb_rd_addr_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_242; // @[Reg.scala 27:20]
  wire [21:0] _T_2862 = _T_2592 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3117 = _T_3116 | _T_2862; // @[Mux.scala 27:72]
  wire  _T_2594 = btb_rd_addr_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_243; // @[Reg.scala 27:20]
  wire [21:0] _T_2863 = _T_2594 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3118 = _T_3117 | _T_2863; // @[Mux.scala 27:72]
  wire  _T_2596 = btb_rd_addr_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_244; // @[Reg.scala 27:20]
  wire [21:0] _T_2864 = _T_2596 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3119 = _T_3118 | _T_2864; // @[Mux.scala 27:72]
  wire  _T_2598 = btb_rd_addr_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_245; // @[Reg.scala 27:20]
  wire [21:0] _T_2865 = _T_2598 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3120 = _T_3119 | _T_2865; // @[Mux.scala 27:72]
  wire  _T_2600 = btb_rd_addr_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_246; // @[Reg.scala 27:20]
  wire [21:0] _T_2866 = _T_2600 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3121 = _T_3120 | _T_2866; // @[Mux.scala 27:72]
  wire  _T_2602 = btb_rd_addr_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_247; // @[Reg.scala 27:20]
  wire [21:0] _T_2867 = _T_2602 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3122 = _T_3121 | _T_2867; // @[Mux.scala 27:72]
  wire  _T_2604 = btb_rd_addr_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_248; // @[Reg.scala 27:20]
  wire [21:0] _T_2868 = _T_2604 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3123 = _T_3122 | _T_2868; // @[Mux.scala 27:72]
  wire  _T_2606 = btb_rd_addr_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_249; // @[Reg.scala 27:20]
  wire [21:0] _T_2869 = _T_2606 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3124 = _T_3123 | _T_2869; // @[Mux.scala 27:72]
  wire  _T_2608 = btb_rd_addr_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_250; // @[Reg.scala 27:20]
  wire [21:0] _T_2870 = _T_2608 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3125 = _T_3124 | _T_2870; // @[Mux.scala 27:72]
  wire  _T_2610 = btb_rd_addr_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_251; // @[Reg.scala 27:20]
  wire [21:0] _T_2871 = _T_2610 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3126 = _T_3125 | _T_2871; // @[Mux.scala 27:72]
  wire  _T_2612 = btb_rd_addr_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_252; // @[Reg.scala 27:20]
  wire [21:0] _T_2872 = _T_2612 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3127 = _T_3126 | _T_2872; // @[Mux.scala 27:72]
  wire  _T_2614 = btb_rd_addr_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_253; // @[Reg.scala 27:20]
  wire [21:0] _T_2873 = _T_2614 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3128 = _T_3127 | _T_2873; // @[Mux.scala 27:72]
  wire  _T_2616 = btb_rd_addr_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_254; // @[Reg.scala 27:20]
  wire [21:0] _T_2874 = _T_2616 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3129 = _T_3128 | _T_2874; // @[Mux.scala 27:72]
  wire  _T_2618 = btb_rd_addr_f == 8'hff; // @[el2_ifu_bp_ctl.scala 368:77]
  reg [21:0] btb_bank0_rd_data_way0_out_255; // @[Reg.scala 27:20]
  wire [21:0] _T_2875 = _T_2618 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_f = _T_3129 | _T_2875; // @[Mux.scala 27:72]
  wire [4:0] _T_25 = io_ifc_fetch_addr_f[13:9] ^ io_ifc_fetch_addr_f[18:14]; // @[el2_lib.scala 177:111]
  wire [4:0] fetch_rd_tag_f = _T_25 ^ io_ifc_fetch_addr_f[23:19]; // @[el2_lib.scala 177:111]
  wire  _T_45 = btb_bank0_rd_data_way0_f[21:17] == fetch_rd_tag_f; // @[el2_ifu_bp_ctl.scala 134:97]
  wire  _T_46 = btb_bank0_rd_data_way0_f[0] & _T_45; // @[el2_ifu_bp_ctl.scala 134:55]
  reg  dec_tlu_way_wb_f; // @[el2_ifu_bp_ctl.scala 126:59]
  wire [6:0] btb_error_addr_wb = io_exu_i0_br_index_r[6:0]; // @[el2_ifu_bp_ctl.scala 93:21]
  wire [7:0] _GEN_1034 = {{1'd0}, btb_error_addr_wb}; // @[el2_ifu_bp_ctl.scala 112:72]
  wire  _T_19 = _GEN_1034 == btb_rd_addr_f; // @[el2_ifu_bp_ctl.scala 112:72]
  wire  branch_error_collision_f = dec_tlu_error_wb & _T_19; // @[el2_ifu_bp_ctl.scala 112:51]
  wire  branch_error_bank_conflict_f = branch_error_collision_f & dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 116:63]
  wire  _T_47 = dec_tlu_way_wb_f & branch_error_bank_conflict_f; // @[el2_ifu_bp_ctl.scala 135:22]
  wire  _T_48 = ~_T_47; // @[el2_ifu_bp_ctl.scala 135:3]
  wire  _T_49 = _T_46 & _T_48; // @[el2_ifu_bp_ctl.scala 134:117]
  wire  _T_50 = _T_49 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 135:54]
  wire  tag_match_way0_f = _T_50 & _T; // @[el2_ifu_bp_ctl.scala 135:75]
  wire  _T_81 = btb_bank0_rd_data_way0_f[3] ^ btb_bank0_rd_data_way0_f[4]; // @[el2_ifu_bp_ctl.scala 147:91]
  wire  _T_82 = tag_match_way0_f & _T_81; // @[el2_ifu_bp_ctl.scala 147:56]
  wire  _T_86 = ~_T_81; // @[el2_ifu_bp_ctl.scala 148:58]
  wire  _T_87 = tag_match_way0_f & _T_86; // @[el2_ifu_bp_ctl.scala 148:56]
  wire [1:0] tag_match_way0_expanded_f = {_T_82,_T_87}; // @[Cat.scala 29:58]
  wire [21:0] _T_126 = tag_match_way0_expanded_f[1] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_0; // @[Reg.scala 27:20]
  wire [21:0] _T_3644 = _T_2108 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_1; // @[Reg.scala 27:20]
  wire [21:0] _T_3645 = _T_2110 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3900 = _T_3644 | _T_3645; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_2; // @[Reg.scala 27:20]
  wire [21:0] _T_3646 = _T_2112 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3901 = _T_3900 | _T_3646; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_3; // @[Reg.scala 27:20]
  wire [21:0] _T_3647 = _T_2114 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3902 = _T_3901 | _T_3647; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_4; // @[Reg.scala 27:20]
  wire [21:0] _T_3648 = _T_2116 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3903 = _T_3902 | _T_3648; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_5; // @[Reg.scala 27:20]
  wire [21:0] _T_3649 = _T_2118 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3904 = _T_3903 | _T_3649; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_6; // @[Reg.scala 27:20]
  wire [21:0] _T_3650 = _T_2120 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3905 = _T_3904 | _T_3650; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_7; // @[Reg.scala 27:20]
  wire [21:0] _T_3651 = _T_2122 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3906 = _T_3905 | _T_3651; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_8; // @[Reg.scala 27:20]
  wire [21:0] _T_3652 = _T_2124 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3907 = _T_3906 | _T_3652; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_9; // @[Reg.scala 27:20]
  wire [21:0] _T_3653 = _T_2126 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3908 = _T_3907 | _T_3653; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_10; // @[Reg.scala 27:20]
  wire [21:0] _T_3654 = _T_2128 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3909 = _T_3908 | _T_3654; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_11; // @[Reg.scala 27:20]
  wire [21:0] _T_3655 = _T_2130 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3910 = _T_3909 | _T_3655; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_12; // @[Reg.scala 27:20]
  wire [21:0] _T_3656 = _T_2132 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3911 = _T_3910 | _T_3656; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_13; // @[Reg.scala 27:20]
  wire [21:0] _T_3657 = _T_2134 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3912 = _T_3911 | _T_3657; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_14; // @[Reg.scala 27:20]
  wire [21:0] _T_3658 = _T_2136 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3913 = _T_3912 | _T_3658; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_15; // @[Reg.scala 27:20]
  wire [21:0] _T_3659 = _T_2138 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3914 = _T_3913 | _T_3659; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_16; // @[Reg.scala 27:20]
  wire [21:0] _T_3660 = _T_2140 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3915 = _T_3914 | _T_3660; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_17; // @[Reg.scala 27:20]
  wire [21:0] _T_3661 = _T_2142 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3916 = _T_3915 | _T_3661; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_18; // @[Reg.scala 27:20]
  wire [21:0] _T_3662 = _T_2144 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3917 = _T_3916 | _T_3662; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_19; // @[Reg.scala 27:20]
  wire [21:0] _T_3663 = _T_2146 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3918 = _T_3917 | _T_3663; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_20; // @[Reg.scala 27:20]
  wire [21:0] _T_3664 = _T_2148 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3919 = _T_3918 | _T_3664; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_21; // @[Reg.scala 27:20]
  wire [21:0] _T_3665 = _T_2150 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3920 = _T_3919 | _T_3665; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_22; // @[Reg.scala 27:20]
  wire [21:0] _T_3666 = _T_2152 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3921 = _T_3920 | _T_3666; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_23; // @[Reg.scala 27:20]
  wire [21:0] _T_3667 = _T_2154 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3922 = _T_3921 | _T_3667; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_24; // @[Reg.scala 27:20]
  wire [21:0] _T_3668 = _T_2156 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3923 = _T_3922 | _T_3668; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_25; // @[Reg.scala 27:20]
  wire [21:0] _T_3669 = _T_2158 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3924 = _T_3923 | _T_3669; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_26; // @[Reg.scala 27:20]
  wire [21:0] _T_3670 = _T_2160 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3925 = _T_3924 | _T_3670; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_27; // @[Reg.scala 27:20]
  wire [21:0] _T_3671 = _T_2162 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3926 = _T_3925 | _T_3671; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_28; // @[Reg.scala 27:20]
  wire [21:0] _T_3672 = _T_2164 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3927 = _T_3926 | _T_3672; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_29; // @[Reg.scala 27:20]
  wire [21:0] _T_3673 = _T_2166 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3928 = _T_3927 | _T_3673; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_30; // @[Reg.scala 27:20]
  wire [21:0] _T_3674 = _T_2168 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3929 = _T_3928 | _T_3674; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_31; // @[Reg.scala 27:20]
  wire [21:0] _T_3675 = _T_2170 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3930 = _T_3929 | _T_3675; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_32; // @[Reg.scala 27:20]
  wire [21:0] _T_3676 = _T_2172 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3931 = _T_3930 | _T_3676; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_33; // @[Reg.scala 27:20]
  wire [21:0] _T_3677 = _T_2174 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3932 = _T_3931 | _T_3677; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_34; // @[Reg.scala 27:20]
  wire [21:0] _T_3678 = _T_2176 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3933 = _T_3932 | _T_3678; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_35; // @[Reg.scala 27:20]
  wire [21:0] _T_3679 = _T_2178 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3934 = _T_3933 | _T_3679; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_36; // @[Reg.scala 27:20]
  wire [21:0] _T_3680 = _T_2180 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3935 = _T_3934 | _T_3680; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_37; // @[Reg.scala 27:20]
  wire [21:0] _T_3681 = _T_2182 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3936 = _T_3935 | _T_3681; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_38; // @[Reg.scala 27:20]
  wire [21:0] _T_3682 = _T_2184 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3937 = _T_3936 | _T_3682; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_39; // @[Reg.scala 27:20]
  wire [21:0] _T_3683 = _T_2186 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3938 = _T_3937 | _T_3683; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_40; // @[Reg.scala 27:20]
  wire [21:0] _T_3684 = _T_2188 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3939 = _T_3938 | _T_3684; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_41; // @[Reg.scala 27:20]
  wire [21:0] _T_3685 = _T_2190 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3940 = _T_3939 | _T_3685; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_42; // @[Reg.scala 27:20]
  wire [21:0] _T_3686 = _T_2192 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3941 = _T_3940 | _T_3686; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_43; // @[Reg.scala 27:20]
  wire [21:0] _T_3687 = _T_2194 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3942 = _T_3941 | _T_3687; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_44; // @[Reg.scala 27:20]
  wire [21:0] _T_3688 = _T_2196 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3943 = _T_3942 | _T_3688; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_45; // @[Reg.scala 27:20]
  wire [21:0] _T_3689 = _T_2198 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3944 = _T_3943 | _T_3689; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_46; // @[Reg.scala 27:20]
  wire [21:0] _T_3690 = _T_2200 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3945 = _T_3944 | _T_3690; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_47; // @[Reg.scala 27:20]
  wire [21:0] _T_3691 = _T_2202 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3946 = _T_3945 | _T_3691; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_48; // @[Reg.scala 27:20]
  wire [21:0] _T_3692 = _T_2204 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3947 = _T_3946 | _T_3692; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_49; // @[Reg.scala 27:20]
  wire [21:0] _T_3693 = _T_2206 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3948 = _T_3947 | _T_3693; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_50; // @[Reg.scala 27:20]
  wire [21:0] _T_3694 = _T_2208 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3949 = _T_3948 | _T_3694; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_51; // @[Reg.scala 27:20]
  wire [21:0] _T_3695 = _T_2210 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3950 = _T_3949 | _T_3695; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_52; // @[Reg.scala 27:20]
  wire [21:0] _T_3696 = _T_2212 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3951 = _T_3950 | _T_3696; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_53; // @[Reg.scala 27:20]
  wire [21:0] _T_3697 = _T_2214 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3952 = _T_3951 | _T_3697; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_54; // @[Reg.scala 27:20]
  wire [21:0] _T_3698 = _T_2216 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3953 = _T_3952 | _T_3698; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_55; // @[Reg.scala 27:20]
  wire [21:0] _T_3699 = _T_2218 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3954 = _T_3953 | _T_3699; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_56; // @[Reg.scala 27:20]
  wire [21:0] _T_3700 = _T_2220 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3955 = _T_3954 | _T_3700; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_57; // @[Reg.scala 27:20]
  wire [21:0] _T_3701 = _T_2222 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3956 = _T_3955 | _T_3701; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_58; // @[Reg.scala 27:20]
  wire [21:0] _T_3702 = _T_2224 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3957 = _T_3956 | _T_3702; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_59; // @[Reg.scala 27:20]
  wire [21:0] _T_3703 = _T_2226 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3958 = _T_3957 | _T_3703; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_60; // @[Reg.scala 27:20]
  wire [21:0] _T_3704 = _T_2228 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3959 = _T_3958 | _T_3704; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_61; // @[Reg.scala 27:20]
  wire [21:0] _T_3705 = _T_2230 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3960 = _T_3959 | _T_3705; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_62; // @[Reg.scala 27:20]
  wire [21:0] _T_3706 = _T_2232 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3961 = _T_3960 | _T_3706; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_63; // @[Reg.scala 27:20]
  wire [21:0] _T_3707 = _T_2234 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3962 = _T_3961 | _T_3707; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_64; // @[Reg.scala 27:20]
  wire [21:0] _T_3708 = _T_2236 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3963 = _T_3962 | _T_3708; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_65; // @[Reg.scala 27:20]
  wire [21:0] _T_3709 = _T_2238 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3964 = _T_3963 | _T_3709; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_66; // @[Reg.scala 27:20]
  wire [21:0] _T_3710 = _T_2240 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3965 = _T_3964 | _T_3710; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_67; // @[Reg.scala 27:20]
  wire [21:0] _T_3711 = _T_2242 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3966 = _T_3965 | _T_3711; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_68; // @[Reg.scala 27:20]
  wire [21:0] _T_3712 = _T_2244 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3967 = _T_3966 | _T_3712; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_69; // @[Reg.scala 27:20]
  wire [21:0] _T_3713 = _T_2246 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3968 = _T_3967 | _T_3713; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_70; // @[Reg.scala 27:20]
  wire [21:0] _T_3714 = _T_2248 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3969 = _T_3968 | _T_3714; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_71; // @[Reg.scala 27:20]
  wire [21:0] _T_3715 = _T_2250 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3970 = _T_3969 | _T_3715; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_72; // @[Reg.scala 27:20]
  wire [21:0] _T_3716 = _T_2252 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3971 = _T_3970 | _T_3716; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_73; // @[Reg.scala 27:20]
  wire [21:0] _T_3717 = _T_2254 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3972 = _T_3971 | _T_3717; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_74; // @[Reg.scala 27:20]
  wire [21:0] _T_3718 = _T_2256 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3973 = _T_3972 | _T_3718; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_75; // @[Reg.scala 27:20]
  wire [21:0] _T_3719 = _T_2258 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3974 = _T_3973 | _T_3719; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_76; // @[Reg.scala 27:20]
  wire [21:0] _T_3720 = _T_2260 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3975 = _T_3974 | _T_3720; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_77; // @[Reg.scala 27:20]
  wire [21:0] _T_3721 = _T_2262 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3976 = _T_3975 | _T_3721; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_78; // @[Reg.scala 27:20]
  wire [21:0] _T_3722 = _T_2264 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3977 = _T_3976 | _T_3722; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_79; // @[Reg.scala 27:20]
  wire [21:0] _T_3723 = _T_2266 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3978 = _T_3977 | _T_3723; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_80; // @[Reg.scala 27:20]
  wire [21:0] _T_3724 = _T_2268 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3979 = _T_3978 | _T_3724; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_81; // @[Reg.scala 27:20]
  wire [21:0] _T_3725 = _T_2270 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3980 = _T_3979 | _T_3725; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_82; // @[Reg.scala 27:20]
  wire [21:0] _T_3726 = _T_2272 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3981 = _T_3980 | _T_3726; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_83; // @[Reg.scala 27:20]
  wire [21:0] _T_3727 = _T_2274 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3982 = _T_3981 | _T_3727; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_84; // @[Reg.scala 27:20]
  wire [21:0] _T_3728 = _T_2276 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3983 = _T_3982 | _T_3728; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_85; // @[Reg.scala 27:20]
  wire [21:0] _T_3729 = _T_2278 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3984 = _T_3983 | _T_3729; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_86; // @[Reg.scala 27:20]
  wire [21:0] _T_3730 = _T_2280 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3985 = _T_3984 | _T_3730; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_87; // @[Reg.scala 27:20]
  wire [21:0] _T_3731 = _T_2282 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3986 = _T_3985 | _T_3731; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_88; // @[Reg.scala 27:20]
  wire [21:0] _T_3732 = _T_2284 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3987 = _T_3986 | _T_3732; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_89; // @[Reg.scala 27:20]
  wire [21:0] _T_3733 = _T_2286 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3988 = _T_3987 | _T_3733; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_90; // @[Reg.scala 27:20]
  wire [21:0] _T_3734 = _T_2288 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3989 = _T_3988 | _T_3734; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_91; // @[Reg.scala 27:20]
  wire [21:0] _T_3735 = _T_2290 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3990 = _T_3989 | _T_3735; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_92; // @[Reg.scala 27:20]
  wire [21:0] _T_3736 = _T_2292 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3991 = _T_3990 | _T_3736; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_93; // @[Reg.scala 27:20]
  wire [21:0] _T_3737 = _T_2294 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3992 = _T_3991 | _T_3737; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_94; // @[Reg.scala 27:20]
  wire [21:0] _T_3738 = _T_2296 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3993 = _T_3992 | _T_3738; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_95; // @[Reg.scala 27:20]
  wire [21:0] _T_3739 = _T_2298 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3994 = _T_3993 | _T_3739; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_96; // @[Reg.scala 27:20]
  wire [21:0] _T_3740 = _T_2300 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3995 = _T_3994 | _T_3740; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_97; // @[Reg.scala 27:20]
  wire [21:0] _T_3741 = _T_2302 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3996 = _T_3995 | _T_3741; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_98; // @[Reg.scala 27:20]
  wire [21:0] _T_3742 = _T_2304 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3997 = _T_3996 | _T_3742; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_99; // @[Reg.scala 27:20]
  wire [21:0] _T_3743 = _T_2306 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3998 = _T_3997 | _T_3743; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_100; // @[Reg.scala 27:20]
  wire [21:0] _T_3744 = _T_2308 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3999 = _T_3998 | _T_3744; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_101; // @[Reg.scala 27:20]
  wire [21:0] _T_3745 = _T_2310 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4000 = _T_3999 | _T_3745; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_102; // @[Reg.scala 27:20]
  wire [21:0] _T_3746 = _T_2312 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4001 = _T_4000 | _T_3746; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_103; // @[Reg.scala 27:20]
  wire [21:0] _T_3747 = _T_2314 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4002 = _T_4001 | _T_3747; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_104; // @[Reg.scala 27:20]
  wire [21:0] _T_3748 = _T_2316 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4003 = _T_4002 | _T_3748; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_105; // @[Reg.scala 27:20]
  wire [21:0] _T_3749 = _T_2318 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4004 = _T_4003 | _T_3749; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_106; // @[Reg.scala 27:20]
  wire [21:0] _T_3750 = _T_2320 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4005 = _T_4004 | _T_3750; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_107; // @[Reg.scala 27:20]
  wire [21:0] _T_3751 = _T_2322 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4006 = _T_4005 | _T_3751; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_108; // @[Reg.scala 27:20]
  wire [21:0] _T_3752 = _T_2324 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4007 = _T_4006 | _T_3752; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_109; // @[Reg.scala 27:20]
  wire [21:0] _T_3753 = _T_2326 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4008 = _T_4007 | _T_3753; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_110; // @[Reg.scala 27:20]
  wire [21:0] _T_3754 = _T_2328 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4009 = _T_4008 | _T_3754; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_111; // @[Reg.scala 27:20]
  wire [21:0] _T_3755 = _T_2330 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4010 = _T_4009 | _T_3755; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_112; // @[Reg.scala 27:20]
  wire [21:0] _T_3756 = _T_2332 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4011 = _T_4010 | _T_3756; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_113; // @[Reg.scala 27:20]
  wire [21:0] _T_3757 = _T_2334 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4012 = _T_4011 | _T_3757; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_114; // @[Reg.scala 27:20]
  wire [21:0] _T_3758 = _T_2336 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4013 = _T_4012 | _T_3758; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_115; // @[Reg.scala 27:20]
  wire [21:0] _T_3759 = _T_2338 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4014 = _T_4013 | _T_3759; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_116; // @[Reg.scala 27:20]
  wire [21:0] _T_3760 = _T_2340 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4015 = _T_4014 | _T_3760; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_117; // @[Reg.scala 27:20]
  wire [21:0] _T_3761 = _T_2342 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4016 = _T_4015 | _T_3761; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_118; // @[Reg.scala 27:20]
  wire [21:0] _T_3762 = _T_2344 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4017 = _T_4016 | _T_3762; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_119; // @[Reg.scala 27:20]
  wire [21:0] _T_3763 = _T_2346 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4018 = _T_4017 | _T_3763; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_120; // @[Reg.scala 27:20]
  wire [21:0] _T_3764 = _T_2348 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4019 = _T_4018 | _T_3764; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_121; // @[Reg.scala 27:20]
  wire [21:0] _T_3765 = _T_2350 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4020 = _T_4019 | _T_3765; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_122; // @[Reg.scala 27:20]
  wire [21:0] _T_3766 = _T_2352 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4021 = _T_4020 | _T_3766; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_123; // @[Reg.scala 27:20]
  wire [21:0] _T_3767 = _T_2354 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4022 = _T_4021 | _T_3767; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_124; // @[Reg.scala 27:20]
  wire [21:0] _T_3768 = _T_2356 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4023 = _T_4022 | _T_3768; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_125; // @[Reg.scala 27:20]
  wire [21:0] _T_3769 = _T_2358 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4024 = _T_4023 | _T_3769; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_126; // @[Reg.scala 27:20]
  wire [21:0] _T_3770 = _T_2360 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4025 = _T_4024 | _T_3770; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_127; // @[Reg.scala 27:20]
  wire [21:0] _T_3771 = _T_2362 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4026 = _T_4025 | _T_3771; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_128; // @[Reg.scala 27:20]
  wire [21:0] _T_3772 = _T_2364 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4027 = _T_4026 | _T_3772; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_129; // @[Reg.scala 27:20]
  wire [21:0] _T_3773 = _T_2366 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4028 = _T_4027 | _T_3773; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_130; // @[Reg.scala 27:20]
  wire [21:0] _T_3774 = _T_2368 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4029 = _T_4028 | _T_3774; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_131; // @[Reg.scala 27:20]
  wire [21:0] _T_3775 = _T_2370 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4030 = _T_4029 | _T_3775; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_132; // @[Reg.scala 27:20]
  wire [21:0] _T_3776 = _T_2372 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4031 = _T_4030 | _T_3776; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_133; // @[Reg.scala 27:20]
  wire [21:0] _T_3777 = _T_2374 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4032 = _T_4031 | _T_3777; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_134; // @[Reg.scala 27:20]
  wire [21:0] _T_3778 = _T_2376 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4033 = _T_4032 | _T_3778; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_135; // @[Reg.scala 27:20]
  wire [21:0] _T_3779 = _T_2378 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4034 = _T_4033 | _T_3779; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_136; // @[Reg.scala 27:20]
  wire [21:0] _T_3780 = _T_2380 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4035 = _T_4034 | _T_3780; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_137; // @[Reg.scala 27:20]
  wire [21:0] _T_3781 = _T_2382 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4036 = _T_4035 | _T_3781; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_138; // @[Reg.scala 27:20]
  wire [21:0] _T_3782 = _T_2384 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4037 = _T_4036 | _T_3782; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_139; // @[Reg.scala 27:20]
  wire [21:0] _T_3783 = _T_2386 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4038 = _T_4037 | _T_3783; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_140; // @[Reg.scala 27:20]
  wire [21:0] _T_3784 = _T_2388 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4039 = _T_4038 | _T_3784; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_141; // @[Reg.scala 27:20]
  wire [21:0] _T_3785 = _T_2390 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4040 = _T_4039 | _T_3785; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_142; // @[Reg.scala 27:20]
  wire [21:0] _T_3786 = _T_2392 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4041 = _T_4040 | _T_3786; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_143; // @[Reg.scala 27:20]
  wire [21:0] _T_3787 = _T_2394 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4042 = _T_4041 | _T_3787; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_144; // @[Reg.scala 27:20]
  wire [21:0] _T_3788 = _T_2396 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4043 = _T_4042 | _T_3788; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_145; // @[Reg.scala 27:20]
  wire [21:0] _T_3789 = _T_2398 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4044 = _T_4043 | _T_3789; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_146; // @[Reg.scala 27:20]
  wire [21:0] _T_3790 = _T_2400 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4045 = _T_4044 | _T_3790; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_147; // @[Reg.scala 27:20]
  wire [21:0] _T_3791 = _T_2402 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4046 = _T_4045 | _T_3791; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_148; // @[Reg.scala 27:20]
  wire [21:0] _T_3792 = _T_2404 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4047 = _T_4046 | _T_3792; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_149; // @[Reg.scala 27:20]
  wire [21:0] _T_3793 = _T_2406 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4048 = _T_4047 | _T_3793; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_150; // @[Reg.scala 27:20]
  wire [21:0] _T_3794 = _T_2408 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4049 = _T_4048 | _T_3794; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_151; // @[Reg.scala 27:20]
  wire [21:0] _T_3795 = _T_2410 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4050 = _T_4049 | _T_3795; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_152; // @[Reg.scala 27:20]
  wire [21:0] _T_3796 = _T_2412 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4051 = _T_4050 | _T_3796; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_153; // @[Reg.scala 27:20]
  wire [21:0] _T_3797 = _T_2414 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4052 = _T_4051 | _T_3797; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_154; // @[Reg.scala 27:20]
  wire [21:0] _T_3798 = _T_2416 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4053 = _T_4052 | _T_3798; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_155; // @[Reg.scala 27:20]
  wire [21:0] _T_3799 = _T_2418 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4054 = _T_4053 | _T_3799; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_156; // @[Reg.scala 27:20]
  wire [21:0] _T_3800 = _T_2420 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4055 = _T_4054 | _T_3800; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_157; // @[Reg.scala 27:20]
  wire [21:0] _T_3801 = _T_2422 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4056 = _T_4055 | _T_3801; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_158; // @[Reg.scala 27:20]
  wire [21:0] _T_3802 = _T_2424 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4057 = _T_4056 | _T_3802; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_159; // @[Reg.scala 27:20]
  wire [21:0] _T_3803 = _T_2426 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4058 = _T_4057 | _T_3803; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_160; // @[Reg.scala 27:20]
  wire [21:0] _T_3804 = _T_2428 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4059 = _T_4058 | _T_3804; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_161; // @[Reg.scala 27:20]
  wire [21:0] _T_3805 = _T_2430 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4060 = _T_4059 | _T_3805; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_162; // @[Reg.scala 27:20]
  wire [21:0] _T_3806 = _T_2432 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4061 = _T_4060 | _T_3806; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_163; // @[Reg.scala 27:20]
  wire [21:0] _T_3807 = _T_2434 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4062 = _T_4061 | _T_3807; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_164; // @[Reg.scala 27:20]
  wire [21:0] _T_3808 = _T_2436 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4063 = _T_4062 | _T_3808; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_165; // @[Reg.scala 27:20]
  wire [21:0] _T_3809 = _T_2438 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4064 = _T_4063 | _T_3809; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_166; // @[Reg.scala 27:20]
  wire [21:0] _T_3810 = _T_2440 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4065 = _T_4064 | _T_3810; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_167; // @[Reg.scala 27:20]
  wire [21:0] _T_3811 = _T_2442 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4066 = _T_4065 | _T_3811; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_168; // @[Reg.scala 27:20]
  wire [21:0] _T_3812 = _T_2444 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4067 = _T_4066 | _T_3812; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_169; // @[Reg.scala 27:20]
  wire [21:0] _T_3813 = _T_2446 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4068 = _T_4067 | _T_3813; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_170; // @[Reg.scala 27:20]
  wire [21:0] _T_3814 = _T_2448 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4069 = _T_4068 | _T_3814; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_171; // @[Reg.scala 27:20]
  wire [21:0] _T_3815 = _T_2450 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4070 = _T_4069 | _T_3815; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_172; // @[Reg.scala 27:20]
  wire [21:0] _T_3816 = _T_2452 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4071 = _T_4070 | _T_3816; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_173; // @[Reg.scala 27:20]
  wire [21:0] _T_3817 = _T_2454 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4072 = _T_4071 | _T_3817; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_174; // @[Reg.scala 27:20]
  wire [21:0] _T_3818 = _T_2456 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4073 = _T_4072 | _T_3818; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_175; // @[Reg.scala 27:20]
  wire [21:0] _T_3819 = _T_2458 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4074 = _T_4073 | _T_3819; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_176; // @[Reg.scala 27:20]
  wire [21:0] _T_3820 = _T_2460 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4075 = _T_4074 | _T_3820; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_177; // @[Reg.scala 27:20]
  wire [21:0] _T_3821 = _T_2462 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4076 = _T_4075 | _T_3821; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_178; // @[Reg.scala 27:20]
  wire [21:0] _T_3822 = _T_2464 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4077 = _T_4076 | _T_3822; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_179; // @[Reg.scala 27:20]
  wire [21:0] _T_3823 = _T_2466 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4078 = _T_4077 | _T_3823; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_180; // @[Reg.scala 27:20]
  wire [21:0] _T_3824 = _T_2468 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4079 = _T_4078 | _T_3824; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_181; // @[Reg.scala 27:20]
  wire [21:0] _T_3825 = _T_2470 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4080 = _T_4079 | _T_3825; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_182; // @[Reg.scala 27:20]
  wire [21:0] _T_3826 = _T_2472 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4081 = _T_4080 | _T_3826; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_183; // @[Reg.scala 27:20]
  wire [21:0] _T_3827 = _T_2474 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4082 = _T_4081 | _T_3827; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_184; // @[Reg.scala 27:20]
  wire [21:0] _T_3828 = _T_2476 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4083 = _T_4082 | _T_3828; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_185; // @[Reg.scala 27:20]
  wire [21:0] _T_3829 = _T_2478 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4084 = _T_4083 | _T_3829; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_186; // @[Reg.scala 27:20]
  wire [21:0] _T_3830 = _T_2480 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4085 = _T_4084 | _T_3830; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_187; // @[Reg.scala 27:20]
  wire [21:0] _T_3831 = _T_2482 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4086 = _T_4085 | _T_3831; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_188; // @[Reg.scala 27:20]
  wire [21:0] _T_3832 = _T_2484 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4087 = _T_4086 | _T_3832; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_189; // @[Reg.scala 27:20]
  wire [21:0] _T_3833 = _T_2486 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4088 = _T_4087 | _T_3833; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_190; // @[Reg.scala 27:20]
  wire [21:0] _T_3834 = _T_2488 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4089 = _T_4088 | _T_3834; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_191; // @[Reg.scala 27:20]
  wire [21:0] _T_3835 = _T_2490 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4090 = _T_4089 | _T_3835; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_192; // @[Reg.scala 27:20]
  wire [21:0] _T_3836 = _T_2492 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4091 = _T_4090 | _T_3836; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_193; // @[Reg.scala 27:20]
  wire [21:0] _T_3837 = _T_2494 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4092 = _T_4091 | _T_3837; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_194; // @[Reg.scala 27:20]
  wire [21:0] _T_3838 = _T_2496 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4093 = _T_4092 | _T_3838; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_195; // @[Reg.scala 27:20]
  wire [21:0] _T_3839 = _T_2498 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4094 = _T_4093 | _T_3839; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_196; // @[Reg.scala 27:20]
  wire [21:0] _T_3840 = _T_2500 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4095 = _T_4094 | _T_3840; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_197; // @[Reg.scala 27:20]
  wire [21:0] _T_3841 = _T_2502 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4096 = _T_4095 | _T_3841; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_198; // @[Reg.scala 27:20]
  wire [21:0] _T_3842 = _T_2504 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4097 = _T_4096 | _T_3842; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_199; // @[Reg.scala 27:20]
  wire [21:0] _T_3843 = _T_2506 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4098 = _T_4097 | _T_3843; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_200; // @[Reg.scala 27:20]
  wire [21:0] _T_3844 = _T_2508 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4099 = _T_4098 | _T_3844; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_201; // @[Reg.scala 27:20]
  wire [21:0] _T_3845 = _T_2510 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4100 = _T_4099 | _T_3845; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_202; // @[Reg.scala 27:20]
  wire [21:0] _T_3846 = _T_2512 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4101 = _T_4100 | _T_3846; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_203; // @[Reg.scala 27:20]
  wire [21:0] _T_3847 = _T_2514 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4102 = _T_4101 | _T_3847; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_204; // @[Reg.scala 27:20]
  wire [21:0] _T_3848 = _T_2516 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4103 = _T_4102 | _T_3848; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_205; // @[Reg.scala 27:20]
  wire [21:0] _T_3849 = _T_2518 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4104 = _T_4103 | _T_3849; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_206; // @[Reg.scala 27:20]
  wire [21:0] _T_3850 = _T_2520 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4105 = _T_4104 | _T_3850; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_207; // @[Reg.scala 27:20]
  wire [21:0] _T_3851 = _T_2522 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4106 = _T_4105 | _T_3851; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_208; // @[Reg.scala 27:20]
  wire [21:0] _T_3852 = _T_2524 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4107 = _T_4106 | _T_3852; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_209; // @[Reg.scala 27:20]
  wire [21:0] _T_3853 = _T_2526 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4108 = _T_4107 | _T_3853; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_210; // @[Reg.scala 27:20]
  wire [21:0] _T_3854 = _T_2528 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4109 = _T_4108 | _T_3854; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_211; // @[Reg.scala 27:20]
  wire [21:0] _T_3855 = _T_2530 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4110 = _T_4109 | _T_3855; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_212; // @[Reg.scala 27:20]
  wire [21:0] _T_3856 = _T_2532 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4111 = _T_4110 | _T_3856; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_213; // @[Reg.scala 27:20]
  wire [21:0] _T_3857 = _T_2534 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4112 = _T_4111 | _T_3857; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_214; // @[Reg.scala 27:20]
  wire [21:0] _T_3858 = _T_2536 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4113 = _T_4112 | _T_3858; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_215; // @[Reg.scala 27:20]
  wire [21:0] _T_3859 = _T_2538 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4114 = _T_4113 | _T_3859; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_216; // @[Reg.scala 27:20]
  wire [21:0] _T_3860 = _T_2540 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4115 = _T_4114 | _T_3860; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_217; // @[Reg.scala 27:20]
  wire [21:0] _T_3861 = _T_2542 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4116 = _T_4115 | _T_3861; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_218; // @[Reg.scala 27:20]
  wire [21:0] _T_3862 = _T_2544 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4117 = _T_4116 | _T_3862; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_219; // @[Reg.scala 27:20]
  wire [21:0] _T_3863 = _T_2546 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4118 = _T_4117 | _T_3863; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_220; // @[Reg.scala 27:20]
  wire [21:0] _T_3864 = _T_2548 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4119 = _T_4118 | _T_3864; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_221; // @[Reg.scala 27:20]
  wire [21:0] _T_3865 = _T_2550 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4120 = _T_4119 | _T_3865; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_222; // @[Reg.scala 27:20]
  wire [21:0] _T_3866 = _T_2552 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4121 = _T_4120 | _T_3866; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_223; // @[Reg.scala 27:20]
  wire [21:0] _T_3867 = _T_2554 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4122 = _T_4121 | _T_3867; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_224; // @[Reg.scala 27:20]
  wire [21:0] _T_3868 = _T_2556 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4123 = _T_4122 | _T_3868; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_225; // @[Reg.scala 27:20]
  wire [21:0] _T_3869 = _T_2558 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4124 = _T_4123 | _T_3869; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_226; // @[Reg.scala 27:20]
  wire [21:0] _T_3870 = _T_2560 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4125 = _T_4124 | _T_3870; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_227; // @[Reg.scala 27:20]
  wire [21:0] _T_3871 = _T_2562 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4126 = _T_4125 | _T_3871; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_228; // @[Reg.scala 27:20]
  wire [21:0] _T_3872 = _T_2564 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4127 = _T_4126 | _T_3872; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_229; // @[Reg.scala 27:20]
  wire [21:0] _T_3873 = _T_2566 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4128 = _T_4127 | _T_3873; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_230; // @[Reg.scala 27:20]
  wire [21:0] _T_3874 = _T_2568 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4129 = _T_4128 | _T_3874; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_231; // @[Reg.scala 27:20]
  wire [21:0] _T_3875 = _T_2570 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4130 = _T_4129 | _T_3875; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_232; // @[Reg.scala 27:20]
  wire [21:0] _T_3876 = _T_2572 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4131 = _T_4130 | _T_3876; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_233; // @[Reg.scala 27:20]
  wire [21:0] _T_3877 = _T_2574 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4132 = _T_4131 | _T_3877; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_234; // @[Reg.scala 27:20]
  wire [21:0] _T_3878 = _T_2576 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4133 = _T_4132 | _T_3878; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_235; // @[Reg.scala 27:20]
  wire [21:0] _T_3879 = _T_2578 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4134 = _T_4133 | _T_3879; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_236; // @[Reg.scala 27:20]
  wire [21:0] _T_3880 = _T_2580 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4135 = _T_4134 | _T_3880; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_237; // @[Reg.scala 27:20]
  wire [21:0] _T_3881 = _T_2582 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4136 = _T_4135 | _T_3881; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_238; // @[Reg.scala 27:20]
  wire [21:0] _T_3882 = _T_2584 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4137 = _T_4136 | _T_3882; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_239; // @[Reg.scala 27:20]
  wire [21:0] _T_3883 = _T_2586 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4138 = _T_4137 | _T_3883; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_240; // @[Reg.scala 27:20]
  wire [21:0] _T_3884 = _T_2588 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4139 = _T_4138 | _T_3884; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_241; // @[Reg.scala 27:20]
  wire [21:0] _T_3885 = _T_2590 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4140 = _T_4139 | _T_3885; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_242; // @[Reg.scala 27:20]
  wire [21:0] _T_3886 = _T_2592 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4141 = _T_4140 | _T_3886; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_243; // @[Reg.scala 27:20]
  wire [21:0] _T_3887 = _T_2594 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4142 = _T_4141 | _T_3887; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_244; // @[Reg.scala 27:20]
  wire [21:0] _T_3888 = _T_2596 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4143 = _T_4142 | _T_3888; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_245; // @[Reg.scala 27:20]
  wire [21:0] _T_3889 = _T_2598 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4144 = _T_4143 | _T_3889; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_246; // @[Reg.scala 27:20]
  wire [21:0] _T_3890 = _T_2600 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4145 = _T_4144 | _T_3890; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_247; // @[Reg.scala 27:20]
  wire [21:0] _T_3891 = _T_2602 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4146 = _T_4145 | _T_3891; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_248; // @[Reg.scala 27:20]
  wire [21:0] _T_3892 = _T_2604 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4147 = _T_4146 | _T_3892; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_249; // @[Reg.scala 27:20]
  wire [21:0] _T_3893 = _T_2606 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4148 = _T_4147 | _T_3893; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_250; // @[Reg.scala 27:20]
  wire [21:0] _T_3894 = _T_2608 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4149 = _T_4148 | _T_3894; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_251; // @[Reg.scala 27:20]
  wire [21:0] _T_3895 = _T_2610 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4150 = _T_4149 | _T_3895; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_252; // @[Reg.scala 27:20]
  wire [21:0] _T_3896 = _T_2612 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4151 = _T_4150 | _T_3896; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_253; // @[Reg.scala 27:20]
  wire [21:0] _T_3897 = _T_2614 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4152 = _T_4151 | _T_3897; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_254; // @[Reg.scala 27:20]
  wire [21:0] _T_3898 = _T_2616 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4153 = _T_4152 | _T_3898; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_255; // @[Reg.scala 27:20]
  wire [21:0] _T_3899 = _T_2618 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_f = _T_4153 | _T_3899; // @[Mux.scala 27:72]
  wire  _T_54 = btb_bank0_rd_data_way1_f[21:17] == fetch_rd_tag_f; // @[el2_ifu_bp_ctl.scala 137:97]
  wire  _T_55 = btb_bank0_rd_data_way1_f[0] & _T_54; // @[el2_ifu_bp_ctl.scala 137:55]
  wire  _T_58 = _T_55 & _T_48; // @[el2_ifu_bp_ctl.scala 137:117]
  wire  _T_59 = _T_58 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 138:54]
  wire  tag_match_way1_f = _T_59 & _T; // @[el2_ifu_bp_ctl.scala 138:75]
  wire  _T_90 = btb_bank0_rd_data_way1_f[3] ^ btb_bank0_rd_data_way1_f[4]; // @[el2_ifu_bp_ctl.scala 150:91]
  wire  _T_91 = tag_match_way1_f & _T_90; // @[el2_ifu_bp_ctl.scala 150:56]
  wire  _T_95 = ~_T_90; // @[el2_ifu_bp_ctl.scala 151:58]
  wire  _T_96 = tag_match_way1_f & _T_95; // @[el2_ifu_bp_ctl.scala 151:56]
  wire [1:0] tag_match_way1_expanded_f = {_T_91,_T_96}; // @[Cat.scala 29:58]
  wire [21:0] _T_127 = tag_match_way1_expanded_f[1] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0o_rd_data_f = _T_126 | _T_127; // @[Mux.scala 27:72]
  wire [21:0] _T_145 = _T_143 ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4156 = btb_rd_addr_p1_f == 8'h0; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4668 = _T_4156 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4158 = btb_rd_addr_p1_f == 8'h1; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4669 = _T_4158 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4924 = _T_4668 | _T_4669; // @[Mux.scala 27:72]
  wire  _T_4160 = btb_rd_addr_p1_f == 8'h2; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4670 = _T_4160 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4925 = _T_4924 | _T_4670; // @[Mux.scala 27:72]
  wire  _T_4162 = btb_rd_addr_p1_f == 8'h3; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4671 = _T_4162 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4926 = _T_4925 | _T_4671; // @[Mux.scala 27:72]
  wire  _T_4164 = btb_rd_addr_p1_f == 8'h4; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4672 = _T_4164 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4927 = _T_4926 | _T_4672; // @[Mux.scala 27:72]
  wire  _T_4166 = btb_rd_addr_p1_f == 8'h5; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4673 = _T_4166 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4928 = _T_4927 | _T_4673; // @[Mux.scala 27:72]
  wire  _T_4168 = btb_rd_addr_p1_f == 8'h6; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4674 = _T_4168 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4929 = _T_4928 | _T_4674; // @[Mux.scala 27:72]
  wire  _T_4170 = btb_rd_addr_p1_f == 8'h7; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4675 = _T_4170 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4930 = _T_4929 | _T_4675; // @[Mux.scala 27:72]
  wire  _T_4172 = btb_rd_addr_p1_f == 8'h8; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4676 = _T_4172 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4931 = _T_4930 | _T_4676; // @[Mux.scala 27:72]
  wire  _T_4174 = btb_rd_addr_p1_f == 8'h9; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4677 = _T_4174 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4932 = _T_4931 | _T_4677; // @[Mux.scala 27:72]
  wire  _T_4176 = btb_rd_addr_p1_f == 8'ha; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4678 = _T_4176 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4933 = _T_4932 | _T_4678; // @[Mux.scala 27:72]
  wire  _T_4178 = btb_rd_addr_p1_f == 8'hb; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4679 = _T_4178 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4934 = _T_4933 | _T_4679; // @[Mux.scala 27:72]
  wire  _T_4180 = btb_rd_addr_p1_f == 8'hc; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4680 = _T_4180 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4935 = _T_4934 | _T_4680; // @[Mux.scala 27:72]
  wire  _T_4182 = btb_rd_addr_p1_f == 8'hd; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4681 = _T_4182 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4936 = _T_4935 | _T_4681; // @[Mux.scala 27:72]
  wire  _T_4184 = btb_rd_addr_p1_f == 8'he; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4682 = _T_4184 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4937 = _T_4936 | _T_4682; // @[Mux.scala 27:72]
  wire  _T_4186 = btb_rd_addr_p1_f == 8'hf; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4683 = _T_4186 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4938 = _T_4937 | _T_4683; // @[Mux.scala 27:72]
  wire  _T_4188 = btb_rd_addr_p1_f == 8'h10; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4684 = _T_4188 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4939 = _T_4938 | _T_4684; // @[Mux.scala 27:72]
  wire  _T_4190 = btb_rd_addr_p1_f == 8'h11; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4685 = _T_4190 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4940 = _T_4939 | _T_4685; // @[Mux.scala 27:72]
  wire  _T_4192 = btb_rd_addr_p1_f == 8'h12; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4686 = _T_4192 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4941 = _T_4940 | _T_4686; // @[Mux.scala 27:72]
  wire  _T_4194 = btb_rd_addr_p1_f == 8'h13; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4687 = _T_4194 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4942 = _T_4941 | _T_4687; // @[Mux.scala 27:72]
  wire  _T_4196 = btb_rd_addr_p1_f == 8'h14; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4688 = _T_4196 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4943 = _T_4942 | _T_4688; // @[Mux.scala 27:72]
  wire  _T_4198 = btb_rd_addr_p1_f == 8'h15; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4689 = _T_4198 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4944 = _T_4943 | _T_4689; // @[Mux.scala 27:72]
  wire  _T_4200 = btb_rd_addr_p1_f == 8'h16; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4690 = _T_4200 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4945 = _T_4944 | _T_4690; // @[Mux.scala 27:72]
  wire  _T_4202 = btb_rd_addr_p1_f == 8'h17; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4691 = _T_4202 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4946 = _T_4945 | _T_4691; // @[Mux.scala 27:72]
  wire  _T_4204 = btb_rd_addr_p1_f == 8'h18; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4692 = _T_4204 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4947 = _T_4946 | _T_4692; // @[Mux.scala 27:72]
  wire  _T_4206 = btb_rd_addr_p1_f == 8'h19; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4693 = _T_4206 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4948 = _T_4947 | _T_4693; // @[Mux.scala 27:72]
  wire  _T_4208 = btb_rd_addr_p1_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4694 = _T_4208 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4949 = _T_4948 | _T_4694; // @[Mux.scala 27:72]
  wire  _T_4210 = btb_rd_addr_p1_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4695 = _T_4210 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4950 = _T_4949 | _T_4695; // @[Mux.scala 27:72]
  wire  _T_4212 = btb_rd_addr_p1_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4696 = _T_4212 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4951 = _T_4950 | _T_4696; // @[Mux.scala 27:72]
  wire  _T_4214 = btb_rd_addr_p1_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4697 = _T_4214 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4952 = _T_4951 | _T_4697; // @[Mux.scala 27:72]
  wire  _T_4216 = btb_rd_addr_p1_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4698 = _T_4216 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4953 = _T_4952 | _T_4698; // @[Mux.scala 27:72]
  wire  _T_4218 = btb_rd_addr_p1_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4699 = _T_4218 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4954 = _T_4953 | _T_4699; // @[Mux.scala 27:72]
  wire  _T_4220 = btb_rd_addr_p1_f == 8'h20; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4700 = _T_4220 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4955 = _T_4954 | _T_4700; // @[Mux.scala 27:72]
  wire  _T_4222 = btb_rd_addr_p1_f == 8'h21; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4701 = _T_4222 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4956 = _T_4955 | _T_4701; // @[Mux.scala 27:72]
  wire  _T_4224 = btb_rd_addr_p1_f == 8'h22; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4702 = _T_4224 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4957 = _T_4956 | _T_4702; // @[Mux.scala 27:72]
  wire  _T_4226 = btb_rd_addr_p1_f == 8'h23; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4703 = _T_4226 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4958 = _T_4957 | _T_4703; // @[Mux.scala 27:72]
  wire  _T_4228 = btb_rd_addr_p1_f == 8'h24; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4704 = _T_4228 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4959 = _T_4958 | _T_4704; // @[Mux.scala 27:72]
  wire  _T_4230 = btb_rd_addr_p1_f == 8'h25; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4705 = _T_4230 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4960 = _T_4959 | _T_4705; // @[Mux.scala 27:72]
  wire  _T_4232 = btb_rd_addr_p1_f == 8'h26; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4706 = _T_4232 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4961 = _T_4960 | _T_4706; // @[Mux.scala 27:72]
  wire  _T_4234 = btb_rd_addr_p1_f == 8'h27; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4707 = _T_4234 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4962 = _T_4961 | _T_4707; // @[Mux.scala 27:72]
  wire  _T_4236 = btb_rd_addr_p1_f == 8'h28; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4708 = _T_4236 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4963 = _T_4962 | _T_4708; // @[Mux.scala 27:72]
  wire  _T_4238 = btb_rd_addr_p1_f == 8'h29; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4709 = _T_4238 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4964 = _T_4963 | _T_4709; // @[Mux.scala 27:72]
  wire  _T_4240 = btb_rd_addr_p1_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4710 = _T_4240 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4965 = _T_4964 | _T_4710; // @[Mux.scala 27:72]
  wire  _T_4242 = btb_rd_addr_p1_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4711 = _T_4242 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4966 = _T_4965 | _T_4711; // @[Mux.scala 27:72]
  wire  _T_4244 = btb_rd_addr_p1_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4712 = _T_4244 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4967 = _T_4966 | _T_4712; // @[Mux.scala 27:72]
  wire  _T_4246 = btb_rd_addr_p1_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4713 = _T_4246 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4968 = _T_4967 | _T_4713; // @[Mux.scala 27:72]
  wire  _T_4248 = btb_rd_addr_p1_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4714 = _T_4248 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4969 = _T_4968 | _T_4714; // @[Mux.scala 27:72]
  wire  _T_4250 = btb_rd_addr_p1_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4715 = _T_4250 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4970 = _T_4969 | _T_4715; // @[Mux.scala 27:72]
  wire  _T_4252 = btb_rd_addr_p1_f == 8'h30; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4716 = _T_4252 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4971 = _T_4970 | _T_4716; // @[Mux.scala 27:72]
  wire  _T_4254 = btb_rd_addr_p1_f == 8'h31; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4717 = _T_4254 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4972 = _T_4971 | _T_4717; // @[Mux.scala 27:72]
  wire  _T_4256 = btb_rd_addr_p1_f == 8'h32; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4718 = _T_4256 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4973 = _T_4972 | _T_4718; // @[Mux.scala 27:72]
  wire  _T_4258 = btb_rd_addr_p1_f == 8'h33; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4719 = _T_4258 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4974 = _T_4973 | _T_4719; // @[Mux.scala 27:72]
  wire  _T_4260 = btb_rd_addr_p1_f == 8'h34; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4720 = _T_4260 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4975 = _T_4974 | _T_4720; // @[Mux.scala 27:72]
  wire  _T_4262 = btb_rd_addr_p1_f == 8'h35; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4721 = _T_4262 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4976 = _T_4975 | _T_4721; // @[Mux.scala 27:72]
  wire  _T_4264 = btb_rd_addr_p1_f == 8'h36; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4722 = _T_4264 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4977 = _T_4976 | _T_4722; // @[Mux.scala 27:72]
  wire  _T_4266 = btb_rd_addr_p1_f == 8'h37; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4723 = _T_4266 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4978 = _T_4977 | _T_4723; // @[Mux.scala 27:72]
  wire  _T_4268 = btb_rd_addr_p1_f == 8'h38; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4724 = _T_4268 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4979 = _T_4978 | _T_4724; // @[Mux.scala 27:72]
  wire  _T_4270 = btb_rd_addr_p1_f == 8'h39; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4725 = _T_4270 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4980 = _T_4979 | _T_4725; // @[Mux.scala 27:72]
  wire  _T_4272 = btb_rd_addr_p1_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4726 = _T_4272 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4981 = _T_4980 | _T_4726; // @[Mux.scala 27:72]
  wire  _T_4274 = btb_rd_addr_p1_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4727 = _T_4274 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4982 = _T_4981 | _T_4727; // @[Mux.scala 27:72]
  wire  _T_4276 = btb_rd_addr_p1_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4728 = _T_4276 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4983 = _T_4982 | _T_4728; // @[Mux.scala 27:72]
  wire  _T_4278 = btb_rd_addr_p1_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4729 = _T_4278 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4984 = _T_4983 | _T_4729; // @[Mux.scala 27:72]
  wire  _T_4280 = btb_rd_addr_p1_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4730 = _T_4280 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4985 = _T_4984 | _T_4730; // @[Mux.scala 27:72]
  wire  _T_4282 = btb_rd_addr_p1_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4731 = _T_4282 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4986 = _T_4985 | _T_4731; // @[Mux.scala 27:72]
  wire  _T_4284 = btb_rd_addr_p1_f == 8'h40; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4732 = _T_4284 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4987 = _T_4986 | _T_4732; // @[Mux.scala 27:72]
  wire  _T_4286 = btb_rd_addr_p1_f == 8'h41; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4733 = _T_4286 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4988 = _T_4987 | _T_4733; // @[Mux.scala 27:72]
  wire  _T_4288 = btb_rd_addr_p1_f == 8'h42; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4734 = _T_4288 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4989 = _T_4988 | _T_4734; // @[Mux.scala 27:72]
  wire  _T_4290 = btb_rd_addr_p1_f == 8'h43; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4735 = _T_4290 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4990 = _T_4989 | _T_4735; // @[Mux.scala 27:72]
  wire  _T_4292 = btb_rd_addr_p1_f == 8'h44; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4736 = _T_4292 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4991 = _T_4990 | _T_4736; // @[Mux.scala 27:72]
  wire  _T_4294 = btb_rd_addr_p1_f == 8'h45; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4737 = _T_4294 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4992 = _T_4991 | _T_4737; // @[Mux.scala 27:72]
  wire  _T_4296 = btb_rd_addr_p1_f == 8'h46; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4738 = _T_4296 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4993 = _T_4992 | _T_4738; // @[Mux.scala 27:72]
  wire  _T_4298 = btb_rd_addr_p1_f == 8'h47; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4739 = _T_4298 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4994 = _T_4993 | _T_4739; // @[Mux.scala 27:72]
  wire  _T_4300 = btb_rd_addr_p1_f == 8'h48; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4740 = _T_4300 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4995 = _T_4994 | _T_4740; // @[Mux.scala 27:72]
  wire  _T_4302 = btb_rd_addr_p1_f == 8'h49; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4741 = _T_4302 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4996 = _T_4995 | _T_4741; // @[Mux.scala 27:72]
  wire  _T_4304 = btb_rd_addr_p1_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4742 = _T_4304 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4997 = _T_4996 | _T_4742; // @[Mux.scala 27:72]
  wire  _T_4306 = btb_rd_addr_p1_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4743 = _T_4306 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4998 = _T_4997 | _T_4743; // @[Mux.scala 27:72]
  wire  _T_4308 = btb_rd_addr_p1_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4744 = _T_4308 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4999 = _T_4998 | _T_4744; // @[Mux.scala 27:72]
  wire  _T_4310 = btb_rd_addr_p1_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4745 = _T_4310 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5000 = _T_4999 | _T_4745; // @[Mux.scala 27:72]
  wire  _T_4312 = btb_rd_addr_p1_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4746 = _T_4312 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5001 = _T_5000 | _T_4746; // @[Mux.scala 27:72]
  wire  _T_4314 = btb_rd_addr_p1_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4747 = _T_4314 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5002 = _T_5001 | _T_4747; // @[Mux.scala 27:72]
  wire  _T_4316 = btb_rd_addr_p1_f == 8'h50; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4748 = _T_4316 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5003 = _T_5002 | _T_4748; // @[Mux.scala 27:72]
  wire  _T_4318 = btb_rd_addr_p1_f == 8'h51; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4749 = _T_4318 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5004 = _T_5003 | _T_4749; // @[Mux.scala 27:72]
  wire  _T_4320 = btb_rd_addr_p1_f == 8'h52; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4750 = _T_4320 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5005 = _T_5004 | _T_4750; // @[Mux.scala 27:72]
  wire  _T_4322 = btb_rd_addr_p1_f == 8'h53; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4751 = _T_4322 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5006 = _T_5005 | _T_4751; // @[Mux.scala 27:72]
  wire  _T_4324 = btb_rd_addr_p1_f == 8'h54; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4752 = _T_4324 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5007 = _T_5006 | _T_4752; // @[Mux.scala 27:72]
  wire  _T_4326 = btb_rd_addr_p1_f == 8'h55; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4753 = _T_4326 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5008 = _T_5007 | _T_4753; // @[Mux.scala 27:72]
  wire  _T_4328 = btb_rd_addr_p1_f == 8'h56; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4754 = _T_4328 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5009 = _T_5008 | _T_4754; // @[Mux.scala 27:72]
  wire  _T_4330 = btb_rd_addr_p1_f == 8'h57; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4755 = _T_4330 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5010 = _T_5009 | _T_4755; // @[Mux.scala 27:72]
  wire  _T_4332 = btb_rd_addr_p1_f == 8'h58; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4756 = _T_4332 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5011 = _T_5010 | _T_4756; // @[Mux.scala 27:72]
  wire  _T_4334 = btb_rd_addr_p1_f == 8'h59; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4757 = _T_4334 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5012 = _T_5011 | _T_4757; // @[Mux.scala 27:72]
  wire  _T_4336 = btb_rd_addr_p1_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4758 = _T_4336 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5013 = _T_5012 | _T_4758; // @[Mux.scala 27:72]
  wire  _T_4338 = btb_rd_addr_p1_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4759 = _T_4338 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5014 = _T_5013 | _T_4759; // @[Mux.scala 27:72]
  wire  _T_4340 = btb_rd_addr_p1_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4760 = _T_4340 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5015 = _T_5014 | _T_4760; // @[Mux.scala 27:72]
  wire  _T_4342 = btb_rd_addr_p1_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4761 = _T_4342 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5016 = _T_5015 | _T_4761; // @[Mux.scala 27:72]
  wire  _T_4344 = btb_rd_addr_p1_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4762 = _T_4344 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5017 = _T_5016 | _T_4762; // @[Mux.scala 27:72]
  wire  _T_4346 = btb_rd_addr_p1_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4763 = _T_4346 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5018 = _T_5017 | _T_4763; // @[Mux.scala 27:72]
  wire  _T_4348 = btb_rd_addr_p1_f == 8'h60; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4764 = _T_4348 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5019 = _T_5018 | _T_4764; // @[Mux.scala 27:72]
  wire  _T_4350 = btb_rd_addr_p1_f == 8'h61; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4765 = _T_4350 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5020 = _T_5019 | _T_4765; // @[Mux.scala 27:72]
  wire  _T_4352 = btb_rd_addr_p1_f == 8'h62; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4766 = _T_4352 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5021 = _T_5020 | _T_4766; // @[Mux.scala 27:72]
  wire  _T_4354 = btb_rd_addr_p1_f == 8'h63; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4767 = _T_4354 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5022 = _T_5021 | _T_4767; // @[Mux.scala 27:72]
  wire  _T_4356 = btb_rd_addr_p1_f == 8'h64; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4768 = _T_4356 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5023 = _T_5022 | _T_4768; // @[Mux.scala 27:72]
  wire  _T_4358 = btb_rd_addr_p1_f == 8'h65; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4769 = _T_4358 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5024 = _T_5023 | _T_4769; // @[Mux.scala 27:72]
  wire  _T_4360 = btb_rd_addr_p1_f == 8'h66; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4770 = _T_4360 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5025 = _T_5024 | _T_4770; // @[Mux.scala 27:72]
  wire  _T_4362 = btb_rd_addr_p1_f == 8'h67; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4771 = _T_4362 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5026 = _T_5025 | _T_4771; // @[Mux.scala 27:72]
  wire  _T_4364 = btb_rd_addr_p1_f == 8'h68; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4772 = _T_4364 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5027 = _T_5026 | _T_4772; // @[Mux.scala 27:72]
  wire  _T_4366 = btb_rd_addr_p1_f == 8'h69; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4773 = _T_4366 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5028 = _T_5027 | _T_4773; // @[Mux.scala 27:72]
  wire  _T_4368 = btb_rd_addr_p1_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4774 = _T_4368 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5029 = _T_5028 | _T_4774; // @[Mux.scala 27:72]
  wire  _T_4370 = btb_rd_addr_p1_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4775 = _T_4370 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5030 = _T_5029 | _T_4775; // @[Mux.scala 27:72]
  wire  _T_4372 = btb_rd_addr_p1_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4776 = _T_4372 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5031 = _T_5030 | _T_4776; // @[Mux.scala 27:72]
  wire  _T_4374 = btb_rd_addr_p1_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4777 = _T_4374 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5032 = _T_5031 | _T_4777; // @[Mux.scala 27:72]
  wire  _T_4376 = btb_rd_addr_p1_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4778 = _T_4376 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5033 = _T_5032 | _T_4778; // @[Mux.scala 27:72]
  wire  _T_4378 = btb_rd_addr_p1_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4779 = _T_4378 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5034 = _T_5033 | _T_4779; // @[Mux.scala 27:72]
  wire  _T_4380 = btb_rd_addr_p1_f == 8'h70; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4780 = _T_4380 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5035 = _T_5034 | _T_4780; // @[Mux.scala 27:72]
  wire  _T_4382 = btb_rd_addr_p1_f == 8'h71; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4781 = _T_4382 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5036 = _T_5035 | _T_4781; // @[Mux.scala 27:72]
  wire  _T_4384 = btb_rd_addr_p1_f == 8'h72; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4782 = _T_4384 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5037 = _T_5036 | _T_4782; // @[Mux.scala 27:72]
  wire  _T_4386 = btb_rd_addr_p1_f == 8'h73; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4783 = _T_4386 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5038 = _T_5037 | _T_4783; // @[Mux.scala 27:72]
  wire  _T_4388 = btb_rd_addr_p1_f == 8'h74; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4784 = _T_4388 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5039 = _T_5038 | _T_4784; // @[Mux.scala 27:72]
  wire  _T_4390 = btb_rd_addr_p1_f == 8'h75; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4785 = _T_4390 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5040 = _T_5039 | _T_4785; // @[Mux.scala 27:72]
  wire  _T_4392 = btb_rd_addr_p1_f == 8'h76; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4786 = _T_4392 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5041 = _T_5040 | _T_4786; // @[Mux.scala 27:72]
  wire  _T_4394 = btb_rd_addr_p1_f == 8'h77; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4787 = _T_4394 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5042 = _T_5041 | _T_4787; // @[Mux.scala 27:72]
  wire  _T_4396 = btb_rd_addr_p1_f == 8'h78; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4788 = _T_4396 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5043 = _T_5042 | _T_4788; // @[Mux.scala 27:72]
  wire  _T_4398 = btb_rd_addr_p1_f == 8'h79; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4789 = _T_4398 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5044 = _T_5043 | _T_4789; // @[Mux.scala 27:72]
  wire  _T_4400 = btb_rd_addr_p1_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4790 = _T_4400 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5045 = _T_5044 | _T_4790; // @[Mux.scala 27:72]
  wire  _T_4402 = btb_rd_addr_p1_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4791 = _T_4402 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5046 = _T_5045 | _T_4791; // @[Mux.scala 27:72]
  wire  _T_4404 = btb_rd_addr_p1_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4792 = _T_4404 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5047 = _T_5046 | _T_4792; // @[Mux.scala 27:72]
  wire  _T_4406 = btb_rd_addr_p1_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4793 = _T_4406 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5048 = _T_5047 | _T_4793; // @[Mux.scala 27:72]
  wire  _T_4408 = btb_rd_addr_p1_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4794 = _T_4408 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5049 = _T_5048 | _T_4794; // @[Mux.scala 27:72]
  wire  _T_4410 = btb_rd_addr_p1_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4795 = _T_4410 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5050 = _T_5049 | _T_4795; // @[Mux.scala 27:72]
  wire  _T_4412 = btb_rd_addr_p1_f == 8'h80; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4796 = _T_4412 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5051 = _T_5050 | _T_4796; // @[Mux.scala 27:72]
  wire  _T_4414 = btb_rd_addr_p1_f == 8'h81; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4797 = _T_4414 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5052 = _T_5051 | _T_4797; // @[Mux.scala 27:72]
  wire  _T_4416 = btb_rd_addr_p1_f == 8'h82; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4798 = _T_4416 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5053 = _T_5052 | _T_4798; // @[Mux.scala 27:72]
  wire  _T_4418 = btb_rd_addr_p1_f == 8'h83; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4799 = _T_4418 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5054 = _T_5053 | _T_4799; // @[Mux.scala 27:72]
  wire  _T_4420 = btb_rd_addr_p1_f == 8'h84; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4800 = _T_4420 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5055 = _T_5054 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4422 = btb_rd_addr_p1_f == 8'h85; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4801 = _T_4422 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5056 = _T_5055 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4424 = btb_rd_addr_p1_f == 8'h86; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4802 = _T_4424 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5057 = _T_5056 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4426 = btb_rd_addr_p1_f == 8'h87; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4803 = _T_4426 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5058 = _T_5057 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4428 = btb_rd_addr_p1_f == 8'h88; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4804 = _T_4428 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5059 = _T_5058 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4430 = btb_rd_addr_p1_f == 8'h89; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4805 = _T_4430 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5060 = _T_5059 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4432 = btb_rd_addr_p1_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4806 = _T_4432 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5061 = _T_5060 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4434 = btb_rd_addr_p1_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4807 = _T_4434 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5062 = _T_5061 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4436 = btb_rd_addr_p1_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4808 = _T_4436 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5063 = _T_5062 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4438 = btb_rd_addr_p1_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4809 = _T_4438 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5064 = _T_5063 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4440 = btb_rd_addr_p1_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4810 = _T_4440 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5065 = _T_5064 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4442 = btb_rd_addr_p1_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4811 = _T_4442 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5066 = _T_5065 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4444 = btb_rd_addr_p1_f == 8'h90; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4812 = _T_4444 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5067 = _T_5066 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4446 = btb_rd_addr_p1_f == 8'h91; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4813 = _T_4446 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5068 = _T_5067 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4448 = btb_rd_addr_p1_f == 8'h92; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4814 = _T_4448 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5069 = _T_5068 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4450 = btb_rd_addr_p1_f == 8'h93; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4815 = _T_4450 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5070 = _T_5069 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4452 = btb_rd_addr_p1_f == 8'h94; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4816 = _T_4452 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5071 = _T_5070 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4454 = btb_rd_addr_p1_f == 8'h95; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4817 = _T_4454 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5072 = _T_5071 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4456 = btb_rd_addr_p1_f == 8'h96; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4818 = _T_4456 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5073 = _T_5072 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4458 = btb_rd_addr_p1_f == 8'h97; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4819 = _T_4458 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5074 = _T_5073 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4460 = btb_rd_addr_p1_f == 8'h98; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4820 = _T_4460 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5075 = _T_5074 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4462 = btb_rd_addr_p1_f == 8'h99; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4821 = _T_4462 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5076 = _T_5075 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4464 = btb_rd_addr_p1_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4822 = _T_4464 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5077 = _T_5076 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4466 = btb_rd_addr_p1_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4823 = _T_4466 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5078 = _T_5077 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4468 = btb_rd_addr_p1_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4824 = _T_4468 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5079 = _T_5078 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4470 = btb_rd_addr_p1_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4825 = _T_4470 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5080 = _T_5079 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4472 = btb_rd_addr_p1_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4826 = _T_4472 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5081 = _T_5080 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4474 = btb_rd_addr_p1_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4827 = _T_4474 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5082 = _T_5081 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4476 = btb_rd_addr_p1_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4828 = _T_4476 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5083 = _T_5082 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4478 = btb_rd_addr_p1_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4829 = _T_4478 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5084 = _T_5083 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4480 = btb_rd_addr_p1_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4830 = _T_4480 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5085 = _T_5084 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4482 = btb_rd_addr_p1_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4831 = _T_4482 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5086 = _T_5085 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4484 = btb_rd_addr_p1_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4832 = _T_4484 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5087 = _T_5086 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4486 = btb_rd_addr_p1_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4833 = _T_4486 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5088 = _T_5087 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4488 = btb_rd_addr_p1_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4834 = _T_4488 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5089 = _T_5088 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4490 = btb_rd_addr_p1_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4835 = _T_4490 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5090 = _T_5089 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4492 = btb_rd_addr_p1_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4836 = _T_4492 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5091 = _T_5090 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4494 = btb_rd_addr_p1_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4837 = _T_4494 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5092 = _T_5091 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4496 = btb_rd_addr_p1_f == 8'haa; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4838 = _T_4496 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5093 = _T_5092 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4498 = btb_rd_addr_p1_f == 8'hab; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4839 = _T_4498 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5094 = _T_5093 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4500 = btb_rd_addr_p1_f == 8'hac; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4840 = _T_4500 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5095 = _T_5094 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4502 = btb_rd_addr_p1_f == 8'had; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4841 = _T_4502 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5096 = _T_5095 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4504 = btb_rd_addr_p1_f == 8'hae; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4842 = _T_4504 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5097 = _T_5096 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4506 = btb_rd_addr_p1_f == 8'haf; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4843 = _T_4506 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5098 = _T_5097 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4508 = btb_rd_addr_p1_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4844 = _T_4508 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5099 = _T_5098 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4510 = btb_rd_addr_p1_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4845 = _T_4510 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5100 = _T_5099 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4512 = btb_rd_addr_p1_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4846 = _T_4512 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5101 = _T_5100 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4514 = btb_rd_addr_p1_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4847 = _T_4514 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5102 = _T_5101 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4516 = btb_rd_addr_p1_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4848 = _T_4516 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5103 = _T_5102 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4518 = btb_rd_addr_p1_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4849 = _T_4518 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5104 = _T_5103 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4520 = btb_rd_addr_p1_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4850 = _T_4520 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5105 = _T_5104 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4522 = btb_rd_addr_p1_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4851 = _T_4522 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5106 = _T_5105 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4524 = btb_rd_addr_p1_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4852 = _T_4524 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5107 = _T_5106 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4526 = btb_rd_addr_p1_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4853 = _T_4526 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5108 = _T_5107 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4528 = btb_rd_addr_p1_f == 8'hba; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4854 = _T_4528 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5109 = _T_5108 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4530 = btb_rd_addr_p1_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4855 = _T_4530 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5110 = _T_5109 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4532 = btb_rd_addr_p1_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4856 = _T_4532 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5111 = _T_5110 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4534 = btb_rd_addr_p1_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4857 = _T_4534 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5112 = _T_5111 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4536 = btb_rd_addr_p1_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4858 = _T_4536 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5113 = _T_5112 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4538 = btb_rd_addr_p1_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4859 = _T_4538 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5114 = _T_5113 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4540 = btb_rd_addr_p1_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4860 = _T_4540 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5115 = _T_5114 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4542 = btb_rd_addr_p1_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4861 = _T_4542 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5116 = _T_5115 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4544 = btb_rd_addr_p1_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4862 = _T_4544 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5117 = _T_5116 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4546 = btb_rd_addr_p1_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4863 = _T_4546 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5118 = _T_5117 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4548 = btb_rd_addr_p1_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4864 = _T_4548 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5119 = _T_5118 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4550 = btb_rd_addr_p1_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4865 = _T_4550 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5120 = _T_5119 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4552 = btb_rd_addr_p1_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4866 = _T_4552 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5121 = _T_5120 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4554 = btb_rd_addr_p1_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4867 = _T_4554 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5122 = _T_5121 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4556 = btb_rd_addr_p1_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4868 = _T_4556 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5123 = _T_5122 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4558 = btb_rd_addr_p1_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4869 = _T_4558 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5124 = _T_5123 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4560 = btb_rd_addr_p1_f == 8'hca; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4870 = _T_4560 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5125 = _T_5124 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4562 = btb_rd_addr_p1_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4871 = _T_4562 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5126 = _T_5125 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4564 = btb_rd_addr_p1_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4872 = _T_4564 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5127 = _T_5126 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4566 = btb_rd_addr_p1_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4873 = _T_4566 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5128 = _T_5127 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4568 = btb_rd_addr_p1_f == 8'hce; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4874 = _T_4568 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5129 = _T_5128 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_4570 = btb_rd_addr_p1_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4875 = _T_4570 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5130 = _T_5129 | _T_4875; // @[Mux.scala 27:72]
  wire  _T_4572 = btb_rd_addr_p1_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4876 = _T_4572 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5131 = _T_5130 | _T_4876; // @[Mux.scala 27:72]
  wire  _T_4574 = btb_rd_addr_p1_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4877 = _T_4574 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5132 = _T_5131 | _T_4877; // @[Mux.scala 27:72]
  wire  _T_4576 = btb_rd_addr_p1_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4878 = _T_4576 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5133 = _T_5132 | _T_4878; // @[Mux.scala 27:72]
  wire  _T_4578 = btb_rd_addr_p1_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4879 = _T_4578 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5134 = _T_5133 | _T_4879; // @[Mux.scala 27:72]
  wire  _T_4580 = btb_rd_addr_p1_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4880 = _T_4580 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5135 = _T_5134 | _T_4880; // @[Mux.scala 27:72]
  wire  _T_4582 = btb_rd_addr_p1_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4881 = _T_4582 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5136 = _T_5135 | _T_4881; // @[Mux.scala 27:72]
  wire  _T_4584 = btb_rd_addr_p1_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4882 = _T_4584 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5137 = _T_5136 | _T_4882; // @[Mux.scala 27:72]
  wire  _T_4586 = btb_rd_addr_p1_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4883 = _T_4586 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5138 = _T_5137 | _T_4883; // @[Mux.scala 27:72]
  wire  _T_4588 = btb_rd_addr_p1_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4884 = _T_4588 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5139 = _T_5138 | _T_4884; // @[Mux.scala 27:72]
  wire  _T_4590 = btb_rd_addr_p1_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4885 = _T_4590 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5140 = _T_5139 | _T_4885; // @[Mux.scala 27:72]
  wire  _T_4592 = btb_rd_addr_p1_f == 8'hda; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4886 = _T_4592 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5141 = _T_5140 | _T_4886; // @[Mux.scala 27:72]
  wire  _T_4594 = btb_rd_addr_p1_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4887 = _T_4594 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5142 = _T_5141 | _T_4887; // @[Mux.scala 27:72]
  wire  _T_4596 = btb_rd_addr_p1_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4888 = _T_4596 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5143 = _T_5142 | _T_4888; // @[Mux.scala 27:72]
  wire  _T_4598 = btb_rd_addr_p1_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4889 = _T_4598 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5144 = _T_5143 | _T_4889; // @[Mux.scala 27:72]
  wire  _T_4600 = btb_rd_addr_p1_f == 8'hde; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4890 = _T_4600 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5145 = _T_5144 | _T_4890; // @[Mux.scala 27:72]
  wire  _T_4602 = btb_rd_addr_p1_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4891 = _T_4602 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5146 = _T_5145 | _T_4891; // @[Mux.scala 27:72]
  wire  _T_4604 = btb_rd_addr_p1_f == 8'he0; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4892 = _T_4604 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5147 = _T_5146 | _T_4892; // @[Mux.scala 27:72]
  wire  _T_4606 = btb_rd_addr_p1_f == 8'he1; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4893 = _T_4606 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5148 = _T_5147 | _T_4893; // @[Mux.scala 27:72]
  wire  _T_4608 = btb_rd_addr_p1_f == 8'he2; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4894 = _T_4608 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5149 = _T_5148 | _T_4894; // @[Mux.scala 27:72]
  wire  _T_4610 = btb_rd_addr_p1_f == 8'he3; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4895 = _T_4610 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5150 = _T_5149 | _T_4895; // @[Mux.scala 27:72]
  wire  _T_4612 = btb_rd_addr_p1_f == 8'he4; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4896 = _T_4612 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5151 = _T_5150 | _T_4896; // @[Mux.scala 27:72]
  wire  _T_4614 = btb_rd_addr_p1_f == 8'he5; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4897 = _T_4614 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5152 = _T_5151 | _T_4897; // @[Mux.scala 27:72]
  wire  _T_4616 = btb_rd_addr_p1_f == 8'he6; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4898 = _T_4616 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5153 = _T_5152 | _T_4898; // @[Mux.scala 27:72]
  wire  _T_4618 = btb_rd_addr_p1_f == 8'he7; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4899 = _T_4618 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5154 = _T_5153 | _T_4899; // @[Mux.scala 27:72]
  wire  _T_4620 = btb_rd_addr_p1_f == 8'he8; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4900 = _T_4620 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5155 = _T_5154 | _T_4900; // @[Mux.scala 27:72]
  wire  _T_4622 = btb_rd_addr_p1_f == 8'he9; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4901 = _T_4622 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5156 = _T_5155 | _T_4901; // @[Mux.scala 27:72]
  wire  _T_4624 = btb_rd_addr_p1_f == 8'hea; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4902 = _T_4624 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5157 = _T_5156 | _T_4902; // @[Mux.scala 27:72]
  wire  _T_4626 = btb_rd_addr_p1_f == 8'heb; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4903 = _T_4626 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5158 = _T_5157 | _T_4903; // @[Mux.scala 27:72]
  wire  _T_4628 = btb_rd_addr_p1_f == 8'hec; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4904 = _T_4628 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5159 = _T_5158 | _T_4904; // @[Mux.scala 27:72]
  wire  _T_4630 = btb_rd_addr_p1_f == 8'hed; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4905 = _T_4630 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5160 = _T_5159 | _T_4905; // @[Mux.scala 27:72]
  wire  _T_4632 = btb_rd_addr_p1_f == 8'hee; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4906 = _T_4632 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5161 = _T_5160 | _T_4906; // @[Mux.scala 27:72]
  wire  _T_4634 = btb_rd_addr_p1_f == 8'hef; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4907 = _T_4634 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5162 = _T_5161 | _T_4907; // @[Mux.scala 27:72]
  wire  _T_4636 = btb_rd_addr_p1_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4908 = _T_4636 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5163 = _T_5162 | _T_4908; // @[Mux.scala 27:72]
  wire  _T_4638 = btb_rd_addr_p1_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4909 = _T_4638 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5164 = _T_5163 | _T_4909; // @[Mux.scala 27:72]
  wire  _T_4640 = btb_rd_addr_p1_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4910 = _T_4640 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5165 = _T_5164 | _T_4910; // @[Mux.scala 27:72]
  wire  _T_4642 = btb_rd_addr_p1_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4911 = _T_4642 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5166 = _T_5165 | _T_4911; // @[Mux.scala 27:72]
  wire  _T_4644 = btb_rd_addr_p1_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4912 = _T_4644 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5167 = _T_5166 | _T_4912; // @[Mux.scala 27:72]
  wire  _T_4646 = btb_rd_addr_p1_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4913 = _T_4646 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5168 = _T_5167 | _T_4913; // @[Mux.scala 27:72]
  wire  _T_4648 = btb_rd_addr_p1_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4914 = _T_4648 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5169 = _T_5168 | _T_4914; // @[Mux.scala 27:72]
  wire  _T_4650 = btb_rd_addr_p1_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4915 = _T_4650 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5170 = _T_5169 | _T_4915; // @[Mux.scala 27:72]
  wire  _T_4652 = btb_rd_addr_p1_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4916 = _T_4652 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5171 = _T_5170 | _T_4916; // @[Mux.scala 27:72]
  wire  _T_4654 = btb_rd_addr_p1_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4917 = _T_4654 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5172 = _T_5171 | _T_4917; // @[Mux.scala 27:72]
  wire  _T_4656 = btb_rd_addr_p1_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4918 = _T_4656 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5173 = _T_5172 | _T_4918; // @[Mux.scala 27:72]
  wire  _T_4658 = btb_rd_addr_p1_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4919 = _T_4658 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5174 = _T_5173 | _T_4919; // @[Mux.scala 27:72]
  wire  _T_4660 = btb_rd_addr_p1_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4920 = _T_4660 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5175 = _T_5174 | _T_4920; // @[Mux.scala 27:72]
  wire  _T_4662 = btb_rd_addr_p1_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4921 = _T_4662 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5176 = _T_5175 | _T_4921; // @[Mux.scala 27:72]
  wire  _T_4664 = btb_rd_addr_p1_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4922 = _T_4664 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5177 = _T_5176 | _T_4922; // @[Mux.scala 27:72]
  wire  _T_4666 = btb_rd_addr_p1_f == 8'hff; // @[el2_ifu_bp_ctl.scala 371:83]
  wire [21:0] _T_4923 = _T_4666 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_p1_f = _T_5177 | _T_4923; // @[Mux.scala 27:72]
  wire [4:0] _T_31 = _T_8[13:9] ^ _T_8[18:14]; // @[el2_lib.scala 177:111]
  wire [4:0] fetch_rd_tag_p1_f = _T_31 ^ _T_8[23:19]; // @[el2_lib.scala 177:111]
  wire  _T_63 = btb_bank0_rd_data_way0_p1_f[21:17] == fetch_rd_tag_p1_f; // @[el2_ifu_bp_ctl.scala 140:106]
  wire  _T_64 = btb_bank0_rd_data_way0_p1_f[0] & _T_63; // @[el2_ifu_bp_ctl.scala 140:61]
  wire  _T_67 = _T_64 & _T_48; // @[el2_ifu_bp_ctl.scala 140:129]
  wire  _T_68 = _T_67 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 141:56]
  wire  tag_match_way0_p1_f = _T_68 & _T; // @[el2_ifu_bp_ctl.scala 141:77]
  wire  _T_99 = btb_bank0_rd_data_way0_p1_f[3] ^ btb_bank0_rd_data_way0_p1_f[4]; // @[el2_ifu_bp_ctl.scala 154:100]
  wire  _T_100 = tag_match_way0_p1_f & _T_99; // @[el2_ifu_bp_ctl.scala 154:62]
  wire  _T_104 = ~_T_99; // @[el2_ifu_bp_ctl.scala 155:64]
  wire  _T_105 = tag_match_way0_p1_f & _T_104; // @[el2_ifu_bp_ctl.scala 155:62]
  wire [1:0] tag_match_way0_expanded_p1_f = {_T_100,_T_105}; // @[Cat.scala 29:58]
  wire [21:0] _T_133 = tag_match_way0_expanded_p1_f[0] ? btb_bank0_rd_data_way0_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5692 = _T_4156 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5693 = _T_4158 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5948 = _T_5692 | _T_5693; // @[Mux.scala 27:72]
  wire [21:0] _T_5694 = _T_4160 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5949 = _T_5948 | _T_5694; // @[Mux.scala 27:72]
  wire [21:0] _T_5695 = _T_4162 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5950 = _T_5949 | _T_5695; // @[Mux.scala 27:72]
  wire [21:0] _T_5696 = _T_4164 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5951 = _T_5950 | _T_5696; // @[Mux.scala 27:72]
  wire [21:0] _T_5697 = _T_4166 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5952 = _T_5951 | _T_5697; // @[Mux.scala 27:72]
  wire [21:0] _T_5698 = _T_4168 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5953 = _T_5952 | _T_5698; // @[Mux.scala 27:72]
  wire [21:0] _T_5699 = _T_4170 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5954 = _T_5953 | _T_5699; // @[Mux.scala 27:72]
  wire [21:0] _T_5700 = _T_4172 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5955 = _T_5954 | _T_5700; // @[Mux.scala 27:72]
  wire [21:0] _T_5701 = _T_4174 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5956 = _T_5955 | _T_5701; // @[Mux.scala 27:72]
  wire [21:0] _T_5702 = _T_4176 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5957 = _T_5956 | _T_5702; // @[Mux.scala 27:72]
  wire [21:0] _T_5703 = _T_4178 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5958 = _T_5957 | _T_5703; // @[Mux.scala 27:72]
  wire [21:0] _T_5704 = _T_4180 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5959 = _T_5958 | _T_5704; // @[Mux.scala 27:72]
  wire [21:0] _T_5705 = _T_4182 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5960 = _T_5959 | _T_5705; // @[Mux.scala 27:72]
  wire [21:0] _T_5706 = _T_4184 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5961 = _T_5960 | _T_5706; // @[Mux.scala 27:72]
  wire [21:0] _T_5707 = _T_4186 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5962 = _T_5961 | _T_5707; // @[Mux.scala 27:72]
  wire [21:0] _T_5708 = _T_4188 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5963 = _T_5962 | _T_5708; // @[Mux.scala 27:72]
  wire [21:0] _T_5709 = _T_4190 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5964 = _T_5963 | _T_5709; // @[Mux.scala 27:72]
  wire [21:0] _T_5710 = _T_4192 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5965 = _T_5964 | _T_5710; // @[Mux.scala 27:72]
  wire [21:0] _T_5711 = _T_4194 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5966 = _T_5965 | _T_5711; // @[Mux.scala 27:72]
  wire [21:0] _T_5712 = _T_4196 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5967 = _T_5966 | _T_5712; // @[Mux.scala 27:72]
  wire [21:0] _T_5713 = _T_4198 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5968 = _T_5967 | _T_5713; // @[Mux.scala 27:72]
  wire [21:0] _T_5714 = _T_4200 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5969 = _T_5968 | _T_5714; // @[Mux.scala 27:72]
  wire [21:0] _T_5715 = _T_4202 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5970 = _T_5969 | _T_5715; // @[Mux.scala 27:72]
  wire [21:0] _T_5716 = _T_4204 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5971 = _T_5970 | _T_5716; // @[Mux.scala 27:72]
  wire [21:0] _T_5717 = _T_4206 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5972 = _T_5971 | _T_5717; // @[Mux.scala 27:72]
  wire [21:0] _T_5718 = _T_4208 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5973 = _T_5972 | _T_5718; // @[Mux.scala 27:72]
  wire [21:0] _T_5719 = _T_4210 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5974 = _T_5973 | _T_5719; // @[Mux.scala 27:72]
  wire [21:0] _T_5720 = _T_4212 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5975 = _T_5974 | _T_5720; // @[Mux.scala 27:72]
  wire [21:0] _T_5721 = _T_4214 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5976 = _T_5975 | _T_5721; // @[Mux.scala 27:72]
  wire [21:0] _T_5722 = _T_4216 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5977 = _T_5976 | _T_5722; // @[Mux.scala 27:72]
  wire [21:0] _T_5723 = _T_4218 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5978 = _T_5977 | _T_5723; // @[Mux.scala 27:72]
  wire [21:0] _T_5724 = _T_4220 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5979 = _T_5978 | _T_5724; // @[Mux.scala 27:72]
  wire [21:0] _T_5725 = _T_4222 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5980 = _T_5979 | _T_5725; // @[Mux.scala 27:72]
  wire [21:0] _T_5726 = _T_4224 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5981 = _T_5980 | _T_5726; // @[Mux.scala 27:72]
  wire [21:0] _T_5727 = _T_4226 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5982 = _T_5981 | _T_5727; // @[Mux.scala 27:72]
  wire [21:0] _T_5728 = _T_4228 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5983 = _T_5982 | _T_5728; // @[Mux.scala 27:72]
  wire [21:0] _T_5729 = _T_4230 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5984 = _T_5983 | _T_5729; // @[Mux.scala 27:72]
  wire [21:0] _T_5730 = _T_4232 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5985 = _T_5984 | _T_5730; // @[Mux.scala 27:72]
  wire [21:0] _T_5731 = _T_4234 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5986 = _T_5985 | _T_5731; // @[Mux.scala 27:72]
  wire [21:0] _T_5732 = _T_4236 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5987 = _T_5986 | _T_5732; // @[Mux.scala 27:72]
  wire [21:0] _T_5733 = _T_4238 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5988 = _T_5987 | _T_5733; // @[Mux.scala 27:72]
  wire [21:0] _T_5734 = _T_4240 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5989 = _T_5988 | _T_5734; // @[Mux.scala 27:72]
  wire [21:0] _T_5735 = _T_4242 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5990 = _T_5989 | _T_5735; // @[Mux.scala 27:72]
  wire [21:0] _T_5736 = _T_4244 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5991 = _T_5990 | _T_5736; // @[Mux.scala 27:72]
  wire [21:0] _T_5737 = _T_4246 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5992 = _T_5991 | _T_5737; // @[Mux.scala 27:72]
  wire [21:0] _T_5738 = _T_4248 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5993 = _T_5992 | _T_5738; // @[Mux.scala 27:72]
  wire [21:0] _T_5739 = _T_4250 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5994 = _T_5993 | _T_5739; // @[Mux.scala 27:72]
  wire [21:0] _T_5740 = _T_4252 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5995 = _T_5994 | _T_5740; // @[Mux.scala 27:72]
  wire [21:0] _T_5741 = _T_4254 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5996 = _T_5995 | _T_5741; // @[Mux.scala 27:72]
  wire [21:0] _T_5742 = _T_4256 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5997 = _T_5996 | _T_5742; // @[Mux.scala 27:72]
  wire [21:0] _T_5743 = _T_4258 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5998 = _T_5997 | _T_5743; // @[Mux.scala 27:72]
  wire [21:0] _T_5744 = _T_4260 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5999 = _T_5998 | _T_5744; // @[Mux.scala 27:72]
  wire [21:0] _T_5745 = _T_4262 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6000 = _T_5999 | _T_5745; // @[Mux.scala 27:72]
  wire [21:0] _T_5746 = _T_4264 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6001 = _T_6000 | _T_5746; // @[Mux.scala 27:72]
  wire [21:0] _T_5747 = _T_4266 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6002 = _T_6001 | _T_5747; // @[Mux.scala 27:72]
  wire [21:0] _T_5748 = _T_4268 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6003 = _T_6002 | _T_5748; // @[Mux.scala 27:72]
  wire [21:0] _T_5749 = _T_4270 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6004 = _T_6003 | _T_5749; // @[Mux.scala 27:72]
  wire [21:0] _T_5750 = _T_4272 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6005 = _T_6004 | _T_5750; // @[Mux.scala 27:72]
  wire [21:0] _T_5751 = _T_4274 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6006 = _T_6005 | _T_5751; // @[Mux.scala 27:72]
  wire [21:0] _T_5752 = _T_4276 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6007 = _T_6006 | _T_5752; // @[Mux.scala 27:72]
  wire [21:0] _T_5753 = _T_4278 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6008 = _T_6007 | _T_5753; // @[Mux.scala 27:72]
  wire [21:0] _T_5754 = _T_4280 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6009 = _T_6008 | _T_5754; // @[Mux.scala 27:72]
  wire [21:0] _T_5755 = _T_4282 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6010 = _T_6009 | _T_5755; // @[Mux.scala 27:72]
  wire [21:0] _T_5756 = _T_4284 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6011 = _T_6010 | _T_5756; // @[Mux.scala 27:72]
  wire [21:0] _T_5757 = _T_4286 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6012 = _T_6011 | _T_5757; // @[Mux.scala 27:72]
  wire [21:0] _T_5758 = _T_4288 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6013 = _T_6012 | _T_5758; // @[Mux.scala 27:72]
  wire [21:0] _T_5759 = _T_4290 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6014 = _T_6013 | _T_5759; // @[Mux.scala 27:72]
  wire [21:0] _T_5760 = _T_4292 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6015 = _T_6014 | _T_5760; // @[Mux.scala 27:72]
  wire [21:0] _T_5761 = _T_4294 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6016 = _T_6015 | _T_5761; // @[Mux.scala 27:72]
  wire [21:0] _T_5762 = _T_4296 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6017 = _T_6016 | _T_5762; // @[Mux.scala 27:72]
  wire [21:0] _T_5763 = _T_4298 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6018 = _T_6017 | _T_5763; // @[Mux.scala 27:72]
  wire [21:0] _T_5764 = _T_4300 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6019 = _T_6018 | _T_5764; // @[Mux.scala 27:72]
  wire [21:0] _T_5765 = _T_4302 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6020 = _T_6019 | _T_5765; // @[Mux.scala 27:72]
  wire [21:0] _T_5766 = _T_4304 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6021 = _T_6020 | _T_5766; // @[Mux.scala 27:72]
  wire [21:0] _T_5767 = _T_4306 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6022 = _T_6021 | _T_5767; // @[Mux.scala 27:72]
  wire [21:0] _T_5768 = _T_4308 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6023 = _T_6022 | _T_5768; // @[Mux.scala 27:72]
  wire [21:0] _T_5769 = _T_4310 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6024 = _T_6023 | _T_5769; // @[Mux.scala 27:72]
  wire [21:0] _T_5770 = _T_4312 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6025 = _T_6024 | _T_5770; // @[Mux.scala 27:72]
  wire [21:0] _T_5771 = _T_4314 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6026 = _T_6025 | _T_5771; // @[Mux.scala 27:72]
  wire [21:0] _T_5772 = _T_4316 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6027 = _T_6026 | _T_5772; // @[Mux.scala 27:72]
  wire [21:0] _T_5773 = _T_4318 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6028 = _T_6027 | _T_5773; // @[Mux.scala 27:72]
  wire [21:0] _T_5774 = _T_4320 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6029 = _T_6028 | _T_5774; // @[Mux.scala 27:72]
  wire [21:0] _T_5775 = _T_4322 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6030 = _T_6029 | _T_5775; // @[Mux.scala 27:72]
  wire [21:0] _T_5776 = _T_4324 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6031 = _T_6030 | _T_5776; // @[Mux.scala 27:72]
  wire [21:0] _T_5777 = _T_4326 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6032 = _T_6031 | _T_5777; // @[Mux.scala 27:72]
  wire [21:0] _T_5778 = _T_4328 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6033 = _T_6032 | _T_5778; // @[Mux.scala 27:72]
  wire [21:0] _T_5779 = _T_4330 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6034 = _T_6033 | _T_5779; // @[Mux.scala 27:72]
  wire [21:0] _T_5780 = _T_4332 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6035 = _T_6034 | _T_5780; // @[Mux.scala 27:72]
  wire [21:0] _T_5781 = _T_4334 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6036 = _T_6035 | _T_5781; // @[Mux.scala 27:72]
  wire [21:0] _T_5782 = _T_4336 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6037 = _T_6036 | _T_5782; // @[Mux.scala 27:72]
  wire [21:0] _T_5783 = _T_4338 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6038 = _T_6037 | _T_5783; // @[Mux.scala 27:72]
  wire [21:0] _T_5784 = _T_4340 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6039 = _T_6038 | _T_5784; // @[Mux.scala 27:72]
  wire [21:0] _T_5785 = _T_4342 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6040 = _T_6039 | _T_5785; // @[Mux.scala 27:72]
  wire [21:0] _T_5786 = _T_4344 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6041 = _T_6040 | _T_5786; // @[Mux.scala 27:72]
  wire [21:0] _T_5787 = _T_4346 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6042 = _T_6041 | _T_5787; // @[Mux.scala 27:72]
  wire [21:0] _T_5788 = _T_4348 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6043 = _T_6042 | _T_5788; // @[Mux.scala 27:72]
  wire [21:0] _T_5789 = _T_4350 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6044 = _T_6043 | _T_5789; // @[Mux.scala 27:72]
  wire [21:0] _T_5790 = _T_4352 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6045 = _T_6044 | _T_5790; // @[Mux.scala 27:72]
  wire [21:0] _T_5791 = _T_4354 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6046 = _T_6045 | _T_5791; // @[Mux.scala 27:72]
  wire [21:0] _T_5792 = _T_4356 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6047 = _T_6046 | _T_5792; // @[Mux.scala 27:72]
  wire [21:0] _T_5793 = _T_4358 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6048 = _T_6047 | _T_5793; // @[Mux.scala 27:72]
  wire [21:0] _T_5794 = _T_4360 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6049 = _T_6048 | _T_5794; // @[Mux.scala 27:72]
  wire [21:0] _T_5795 = _T_4362 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6050 = _T_6049 | _T_5795; // @[Mux.scala 27:72]
  wire [21:0] _T_5796 = _T_4364 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6051 = _T_6050 | _T_5796; // @[Mux.scala 27:72]
  wire [21:0] _T_5797 = _T_4366 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6052 = _T_6051 | _T_5797; // @[Mux.scala 27:72]
  wire [21:0] _T_5798 = _T_4368 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6053 = _T_6052 | _T_5798; // @[Mux.scala 27:72]
  wire [21:0] _T_5799 = _T_4370 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6054 = _T_6053 | _T_5799; // @[Mux.scala 27:72]
  wire [21:0] _T_5800 = _T_4372 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6055 = _T_6054 | _T_5800; // @[Mux.scala 27:72]
  wire [21:0] _T_5801 = _T_4374 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6056 = _T_6055 | _T_5801; // @[Mux.scala 27:72]
  wire [21:0] _T_5802 = _T_4376 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6057 = _T_6056 | _T_5802; // @[Mux.scala 27:72]
  wire [21:0] _T_5803 = _T_4378 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6058 = _T_6057 | _T_5803; // @[Mux.scala 27:72]
  wire [21:0] _T_5804 = _T_4380 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6059 = _T_6058 | _T_5804; // @[Mux.scala 27:72]
  wire [21:0] _T_5805 = _T_4382 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6060 = _T_6059 | _T_5805; // @[Mux.scala 27:72]
  wire [21:0] _T_5806 = _T_4384 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6061 = _T_6060 | _T_5806; // @[Mux.scala 27:72]
  wire [21:0] _T_5807 = _T_4386 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6062 = _T_6061 | _T_5807; // @[Mux.scala 27:72]
  wire [21:0] _T_5808 = _T_4388 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6063 = _T_6062 | _T_5808; // @[Mux.scala 27:72]
  wire [21:0] _T_5809 = _T_4390 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6064 = _T_6063 | _T_5809; // @[Mux.scala 27:72]
  wire [21:0] _T_5810 = _T_4392 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6065 = _T_6064 | _T_5810; // @[Mux.scala 27:72]
  wire [21:0] _T_5811 = _T_4394 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6066 = _T_6065 | _T_5811; // @[Mux.scala 27:72]
  wire [21:0] _T_5812 = _T_4396 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6067 = _T_6066 | _T_5812; // @[Mux.scala 27:72]
  wire [21:0] _T_5813 = _T_4398 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6068 = _T_6067 | _T_5813; // @[Mux.scala 27:72]
  wire [21:0] _T_5814 = _T_4400 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6069 = _T_6068 | _T_5814; // @[Mux.scala 27:72]
  wire [21:0] _T_5815 = _T_4402 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6070 = _T_6069 | _T_5815; // @[Mux.scala 27:72]
  wire [21:0] _T_5816 = _T_4404 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6071 = _T_6070 | _T_5816; // @[Mux.scala 27:72]
  wire [21:0] _T_5817 = _T_4406 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6072 = _T_6071 | _T_5817; // @[Mux.scala 27:72]
  wire [21:0] _T_5818 = _T_4408 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6073 = _T_6072 | _T_5818; // @[Mux.scala 27:72]
  wire [21:0] _T_5819 = _T_4410 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6074 = _T_6073 | _T_5819; // @[Mux.scala 27:72]
  wire [21:0] _T_5820 = _T_4412 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6075 = _T_6074 | _T_5820; // @[Mux.scala 27:72]
  wire [21:0] _T_5821 = _T_4414 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6076 = _T_6075 | _T_5821; // @[Mux.scala 27:72]
  wire [21:0] _T_5822 = _T_4416 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6077 = _T_6076 | _T_5822; // @[Mux.scala 27:72]
  wire [21:0] _T_5823 = _T_4418 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6078 = _T_6077 | _T_5823; // @[Mux.scala 27:72]
  wire [21:0] _T_5824 = _T_4420 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6079 = _T_6078 | _T_5824; // @[Mux.scala 27:72]
  wire [21:0] _T_5825 = _T_4422 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6080 = _T_6079 | _T_5825; // @[Mux.scala 27:72]
  wire [21:0] _T_5826 = _T_4424 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6081 = _T_6080 | _T_5826; // @[Mux.scala 27:72]
  wire [21:0] _T_5827 = _T_4426 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6082 = _T_6081 | _T_5827; // @[Mux.scala 27:72]
  wire [21:0] _T_5828 = _T_4428 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6083 = _T_6082 | _T_5828; // @[Mux.scala 27:72]
  wire [21:0] _T_5829 = _T_4430 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6084 = _T_6083 | _T_5829; // @[Mux.scala 27:72]
  wire [21:0] _T_5830 = _T_4432 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6085 = _T_6084 | _T_5830; // @[Mux.scala 27:72]
  wire [21:0] _T_5831 = _T_4434 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6086 = _T_6085 | _T_5831; // @[Mux.scala 27:72]
  wire [21:0] _T_5832 = _T_4436 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6087 = _T_6086 | _T_5832; // @[Mux.scala 27:72]
  wire [21:0] _T_5833 = _T_4438 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6088 = _T_6087 | _T_5833; // @[Mux.scala 27:72]
  wire [21:0] _T_5834 = _T_4440 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6089 = _T_6088 | _T_5834; // @[Mux.scala 27:72]
  wire [21:0] _T_5835 = _T_4442 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6090 = _T_6089 | _T_5835; // @[Mux.scala 27:72]
  wire [21:0] _T_5836 = _T_4444 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6091 = _T_6090 | _T_5836; // @[Mux.scala 27:72]
  wire [21:0] _T_5837 = _T_4446 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6092 = _T_6091 | _T_5837; // @[Mux.scala 27:72]
  wire [21:0] _T_5838 = _T_4448 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6093 = _T_6092 | _T_5838; // @[Mux.scala 27:72]
  wire [21:0] _T_5839 = _T_4450 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6094 = _T_6093 | _T_5839; // @[Mux.scala 27:72]
  wire [21:0] _T_5840 = _T_4452 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6095 = _T_6094 | _T_5840; // @[Mux.scala 27:72]
  wire [21:0] _T_5841 = _T_4454 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6096 = _T_6095 | _T_5841; // @[Mux.scala 27:72]
  wire [21:0] _T_5842 = _T_4456 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6097 = _T_6096 | _T_5842; // @[Mux.scala 27:72]
  wire [21:0] _T_5843 = _T_4458 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6098 = _T_6097 | _T_5843; // @[Mux.scala 27:72]
  wire [21:0] _T_5844 = _T_4460 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6099 = _T_6098 | _T_5844; // @[Mux.scala 27:72]
  wire [21:0] _T_5845 = _T_4462 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6100 = _T_6099 | _T_5845; // @[Mux.scala 27:72]
  wire [21:0] _T_5846 = _T_4464 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6101 = _T_6100 | _T_5846; // @[Mux.scala 27:72]
  wire [21:0] _T_5847 = _T_4466 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6102 = _T_6101 | _T_5847; // @[Mux.scala 27:72]
  wire [21:0] _T_5848 = _T_4468 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6103 = _T_6102 | _T_5848; // @[Mux.scala 27:72]
  wire [21:0] _T_5849 = _T_4470 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6104 = _T_6103 | _T_5849; // @[Mux.scala 27:72]
  wire [21:0] _T_5850 = _T_4472 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6105 = _T_6104 | _T_5850; // @[Mux.scala 27:72]
  wire [21:0] _T_5851 = _T_4474 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6106 = _T_6105 | _T_5851; // @[Mux.scala 27:72]
  wire [21:0] _T_5852 = _T_4476 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6107 = _T_6106 | _T_5852; // @[Mux.scala 27:72]
  wire [21:0] _T_5853 = _T_4478 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6108 = _T_6107 | _T_5853; // @[Mux.scala 27:72]
  wire [21:0] _T_5854 = _T_4480 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6109 = _T_6108 | _T_5854; // @[Mux.scala 27:72]
  wire [21:0] _T_5855 = _T_4482 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6110 = _T_6109 | _T_5855; // @[Mux.scala 27:72]
  wire [21:0] _T_5856 = _T_4484 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6111 = _T_6110 | _T_5856; // @[Mux.scala 27:72]
  wire [21:0] _T_5857 = _T_4486 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6112 = _T_6111 | _T_5857; // @[Mux.scala 27:72]
  wire [21:0] _T_5858 = _T_4488 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6113 = _T_6112 | _T_5858; // @[Mux.scala 27:72]
  wire [21:0] _T_5859 = _T_4490 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6114 = _T_6113 | _T_5859; // @[Mux.scala 27:72]
  wire [21:0] _T_5860 = _T_4492 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6115 = _T_6114 | _T_5860; // @[Mux.scala 27:72]
  wire [21:0] _T_5861 = _T_4494 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6116 = _T_6115 | _T_5861; // @[Mux.scala 27:72]
  wire [21:0] _T_5862 = _T_4496 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6117 = _T_6116 | _T_5862; // @[Mux.scala 27:72]
  wire [21:0] _T_5863 = _T_4498 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6118 = _T_6117 | _T_5863; // @[Mux.scala 27:72]
  wire [21:0] _T_5864 = _T_4500 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6119 = _T_6118 | _T_5864; // @[Mux.scala 27:72]
  wire [21:0] _T_5865 = _T_4502 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6120 = _T_6119 | _T_5865; // @[Mux.scala 27:72]
  wire [21:0] _T_5866 = _T_4504 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6121 = _T_6120 | _T_5866; // @[Mux.scala 27:72]
  wire [21:0] _T_5867 = _T_4506 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6122 = _T_6121 | _T_5867; // @[Mux.scala 27:72]
  wire [21:0] _T_5868 = _T_4508 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6123 = _T_6122 | _T_5868; // @[Mux.scala 27:72]
  wire [21:0] _T_5869 = _T_4510 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6124 = _T_6123 | _T_5869; // @[Mux.scala 27:72]
  wire [21:0] _T_5870 = _T_4512 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6125 = _T_6124 | _T_5870; // @[Mux.scala 27:72]
  wire [21:0] _T_5871 = _T_4514 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6126 = _T_6125 | _T_5871; // @[Mux.scala 27:72]
  wire [21:0] _T_5872 = _T_4516 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6127 = _T_6126 | _T_5872; // @[Mux.scala 27:72]
  wire [21:0] _T_5873 = _T_4518 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6128 = _T_6127 | _T_5873; // @[Mux.scala 27:72]
  wire [21:0] _T_5874 = _T_4520 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6129 = _T_6128 | _T_5874; // @[Mux.scala 27:72]
  wire [21:0] _T_5875 = _T_4522 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6130 = _T_6129 | _T_5875; // @[Mux.scala 27:72]
  wire [21:0] _T_5876 = _T_4524 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6131 = _T_6130 | _T_5876; // @[Mux.scala 27:72]
  wire [21:0] _T_5877 = _T_4526 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6132 = _T_6131 | _T_5877; // @[Mux.scala 27:72]
  wire [21:0] _T_5878 = _T_4528 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6133 = _T_6132 | _T_5878; // @[Mux.scala 27:72]
  wire [21:0] _T_5879 = _T_4530 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6134 = _T_6133 | _T_5879; // @[Mux.scala 27:72]
  wire [21:0] _T_5880 = _T_4532 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6135 = _T_6134 | _T_5880; // @[Mux.scala 27:72]
  wire [21:0] _T_5881 = _T_4534 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6136 = _T_6135 | _T_5881; // @[Mux.scala 27:72]
  wire [21:0] _T_5882 = _T_4536 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6137 = _T_6136 | _T_5882; // @[Mux.scala 27:72]
  wire [21:0] _T_5883 = _T_4538 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6138 = _T_6137 | _T_5883; // @[Mux.scala 27:72]
  wire [21:0] _T_5884 = _T_4540 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6139 = _T_6138 | _T_5884; // @[Mux.scala 27:72]
  wire [21:0] _T_5885 = _T_4542 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6140 = _T_6139 | _T_5885; // @[Mux.scala 27:72]
  wire [21:0] _T_5886 = _T_4544 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6141 = _T_6140 | _T_5886; // @[Mux.scala 27:72]
  wire [21:0] _T_5887 = _T_4546 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6142 = _T_6141 | _T_5887; // @[Mux.scala 27:72]
  wire [21:0] _T_5888 = _T_4548 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6143 = _T_6142 | _T_5888; // @[Mux.scala 27:72]
  wire [21:0] _T_5889 = _T_4550 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6144 = _T_6143 | _T_5889; // @[Mux.scala 27:72]
  wire [21:0] _T_5890 = _T_4552 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6145 = _T_6144 | _T_5890; // @[Mux.scala 27:72]
  wire [21:0] _T_5891 = _T_4554 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6146 = _T_6145 | _T_5891; // @[Mux.scala 27:72]
  wire [21:0] _T_5892 = _T_4556 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6147 = _T_6146 | _T_5892; // @[Mux.scala 27:72]
  wire [21:0] _T_5893 = _T_4558 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6148 = _T_6147 | _T_5893; // @[Mux.scala 27:72]
  wire [21:0] _T_5894 = _T_4560 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6149 = _T_6148 | _T_5894; // @[Mux.scala 27:72]
  wire [21:0] _T_5895 = _T_4562 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6150 = _T_6149 | _T_5895; // @[Mux.scala 27:72]
  wire [21:0] _T_5896 = _T_4564 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6151 = _T_6150 | _T_5896; // @[Mux.scala 27:72]
  wire [21:0] _T_5897 = _T_4566 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6152 = _T_6151 | _T_5897; // @[Mux.scala 27:72]
  wire [21:0] _T_5898 = _T_4568 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6153 = _T_6152 | _T_5898; // @[Mux.scala 27:72]
  wire [21:0] _T_5899 = _T_4570 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6154 = _T_6153 | _T_5899; // @[Mux.scala 27:72]
  wire [21:0] _T_5900 = _T_4572 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6155 = _T_6154 | _T_5900; // @[Mux.scala 27:72]
  wire [21:0] _T_5901 = _T_4574 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6156 = _T_6155 | _T_5901; // @[Mux.scala 27:72]
  wire [21:0] _T_5902 = _T_4576 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6157 = _T_6156 | _T_5902; // @[Mux.scala 27:72]
  wire [21:0] _T_5903 = _T_4578 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6158 = _T_6157 | _T_5903; // @[Mux.scala 27:72]
  wire [21:0] _T_5904 = _T_4580 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6159 = _T_6158 | _T_5904; // @[Mux.scala 27:72]
  wire [21:0] _T_5905 = _T_4582 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6160 = _T_6159 | _T_5905; // @[Mux.scala 27:72]
  wire [21:0] _T_5906 = _T_4584 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6161 = _T_6160 | _T_5906; // @[Mux.scala 27:72]
  wire [21:0] _T_5907 = _T_4586 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6162 = _T_6161 | _T_5907; // @[Mux.scala 27:72]
  wire [21:0] _T_5908 = _T_4588 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6163 = _T_6162 | _T_5908; // @[Mux.scala 27:72]
  wire [21:0] _T_5909 = _T_4590 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6164 = _T_6163 | _T_5909; // @[Mux.scala 27:72]
  wire [21:0] _T_5910 = _T_4592 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6165 = _T_6164 | _T_5910; // @[Mux.scala 27:72]
  wire [21:0] _T_5911 = _T_4594 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6166 = _T_6165 | _T_5911; // @[Mux.scala 27:72]
  wire [21:0] _T_5912 = _T_4596 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6167 = _T_6166 | _T_5912; // @[Mux.scala 27:72]
  wire [21:0] _T_5913 = _T_4598 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6168 = _T_6167 | _T_5913; // @[Mux.scala 27:72]
  wire [21:0] _T_5914 = _T_4600 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6169 = _T_6168 | _T_5914; // @[Mux.scala 27:72]
  wire [21:0] _T_5915 = _T_4602 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6170 = _T_6169 | _T_5915; // @[Mux.scala 27:72]
  wire [21:0] _T_5916 = _T_4604 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6171 = _T_6170 | _T_5916; // @[Mux.scala 27:72]
  wire [21:0] _T_5917 = _T_4606 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6172 = _T_6171 | _T_5917; // @[Mux.scala 27:72]
  wire [21:0] _T_5918 = _T_4608 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6173 = _T_6172 | _T_5918; // @[Mux.scala 27:72]
  wire [21:0] _T_5919 = _T_4610 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6174 = _T_6173 | _T_5919; // @[Mux.scala 27:72]
  wire [21:0] _T_5920 = _T_4612 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6175 = _T_6174 | _T_5920; // @[Mux.scala 27:72]
  wire [21:0] _T_5921 = _T_4614 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6176 = _T_6175 | _T_5921; // @[Mux.scala 27:72]
  wire [21:0] _T_5922 = _T_4616 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6177 = _T_6176 | _T_5922; // @[Mux.scala 27:72]
  wire [21:0] _T_5923 = _T_4618 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6178 = _T_6177 | _T_5923; // @[Mux.scala 27:72]
  wire [21:0] _T_5924 = _T_4620 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6179 = _T_6178 | _T_5924; // @[Mux.scala 27:72]
  wire [21:0] _T_5925 = _T_4622 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6180 = _T_6179 | _T_5925; // @[Mux.scala 27:72]
  wire [21:0] _T_5926 = _T_4624 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6181 = _T_6180 | _T_5926; // @[Mux.scala 27:72]
  wire [21:0] _T_5927 = _T_4626 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6182 = _T_6181 | _T_5927; // @[Mux.scala 27:72]
  wire [21:0] _T_5928 = _T_4628 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6183 = _T_6182 | _T_5928; // @[Mux.scala 27:72]
  wire [21:0] _T_5929 = _T_4630 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6184 = _T_6183 | _T_5929; // @[Mux.scala 27:72]
  wire [21:0] _T_5930 = _T_4632 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6185 = _T_6184 | _T_5930; // @[Mux.scala 27:72]
  wire [21:0] _T_5931 = _T_4634 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6186 = _T_6185 | _T_5931; // @[Mux.scala 27:72]
  wire [21:0] _T_5932 = _T_4636 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6187 = _T_6186 | _T_5932; // @[Mux.scala 27:72]
  wire [21:0] _T_5933 = _T_4638 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6188 = _T_6187 | _T_5933; // @[Mux.scala 27:72]
  wire [21:0] _T_5934 = _T_4640 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6189 = _T_6188 | _T_5934; // @[Mux.scala 27:72]
  wire [21:0] _T_5935 = _T_4642 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6190 = _T_6189 | _T_5935; // @[Mux.scala 27:72]
  wire [21:0] _T_5936 = _T_4644 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6191 = _T_6190 | _T_5936; // @[Mux.scala 27:72]
  wire [21:0] _T_5937 = _T_4646 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6192 = _T_6191 | _T_5937; // @[Mux.scala 27:72]
  wire [21:0] _T_5938 = _T_4648 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6193 = _T_6192 | _T_5938; // @[Mux.scala 27:72]
  wire [21:0] _T_5939 = _T_4650 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6194 = _T_6193 | _T_5939; // @[Mux.scala 27:72]
  wire [21:0] _T_5940 = _T_4652 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6195 = _T_6194 | _T_5940; // @[Mux.scala 27:72]
  wire [21:0] _T_5941 = _T_4654 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6196 = _T_6195 | _T_5941; // @[Mux.scala 27:72]
  wire [21:0] _T_5942 = _T_4656 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6197 = _T_6196 | _T_5942; // @[Mux.scala 27:72]
  wire [21:0] _T_5943 = _T_4658 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6198 = _T_6197 | _T_5943; // @[Mux.scala 27:72]
  wire [21:0] _T_5944 = _T_4660 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6199 = _T_6198 | _T_5944; // @[Mux.scala 27:72]
  wire [21:0] _T_5945 = _T_4662 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6200 = _T_6199 | _T_5945; // @[Mux.scala 27:72]
  wire [21:0] _T_5946 = _T_4664 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6201 = _T_6200 | _T_5946; // @[Mux.scala 27:72]
  wire [21:0] _T_5947 = _T_4666 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_p1_f = _T_6201 | _T_5947; // @[Mux.scala 27:72]
  wire  _T_72 = btb_bank0_rd_data_way1_p1_f[21:17] == fetch_rd_tag_p1_f; // @[el2_ifu_bp_ctl.scala 143:106]
  wire  _T_73 = btb_bank0_rd_data_way1_p1_f[0] & _T_72; // @[el2_ifu_bp_ctl.scala 143:61]
  wire  _T_76 = _T_73 & _T_48; // @[el2_ifu_bp_ctl.scala 143:129]
  wire  _T_77 = _T_76 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 144:56]
  wire  tag_match_way1_p1_f = _T_77 & _T; // @[el2_ifu_bp_ctl.scala 144:77]
  wire  _T_108 = btb_bank0_rd_data_way1_p1_f[3] ^ btb_bank0_rd_data_way1_p1_f[4]; // @[el2_ifu_bp_ctl.scala 157:100]
  wire  _T_109 = tag_match_way1_p1_f & _T_108; // @[el2_ifu_bp_ctl.scala 157:62]
  wire  _T_113 = ~_T_108; // @[el2_ifu_bp_ctl.scala 158:64]
  wire  _T_114 = tag_match_way1_p1_f & _T_113; // @[el2_ifu_bp_ctl.scala 158:62]
  wire [1:0] tag_match_way1_expanded_p1_f = {_T_109,_T_114}; // @[Cat.scala 29:58]
  wire [21:0] _T_134 = tag_match_way1_expanded_p1_f[0] ? btb_bank0_rd_data_way1_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_p1_f = _T_133 | _T_134; // @[Mux.scala 27:72]
  wire [21:0] _T_146 = io_ifc_fetch_addr_f[0] ? btb_bank0e_rd_data_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank1_rd_data_f = _T_145 | _T_146; // @[Mux.scala 27:72]
  wire  _T_241 = btb_vbank1_rd_data_f[2] | btb_vbank1_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 235:59]
  wire [21:0] _T_119 = tag_match_way0_expanded_f[0] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_120 = tag_match_way1_expanded_f[0] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_f = _T_119 | _T_120; // @[Mux.scala 27:72]
  wire [21:0] _T_139 = _T_143 ? btb_bank0e_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_140 = io_ifc_fetch_addr_f[0] ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank0_rd_data_f = _T_139 | _T_140; // @[Mux.scala 27:72]
  wire  _T_244 = btb_vbank0_rd_data_f[2] | btb_vbank0_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 236:59]
  wire [1:0] bht_force_taken_f = {_T_241,_T_244}; // @[Cat.scala 29:58]
  wire [9:0] _T_566 = {btb_rd_addr_f,2'h0}; // @[Cat.scala 29:58]
  reg [7:0] fghr; // @[el2_ifu_bp_ctl.scala 283:44]
  wire [7:0] bht_rd_addr_hashed_f = _T_566[9:2] ^ fghr; // @[el2_lib.scala 191:35]
  wire  _T_21597 = bht_rd_addr_hashed_f == 8'h0; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_0; // @[Reg.scala 27:20]
  wire [1:0] _T_22364 = _T_21597 ? bht_bank_rd_data_out_1_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_21600 = bht_rd_addr_hashed_f == 8'h1; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_1; // @[Reg.scala 27:20]
  wire [1:0] _T_22365 = _T_21600 ? bht_bank_rd_data_out_1_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22620 = _T_22364 | _T_22365; // @[Mux.scala 27:72]
  wire  _T_21603 = bht_rd_addr_hashed_f == 8'h2; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_2; // @[Reg.scala 27:20]
  wire [1:0] _T_22366 = _T_21603 ? bht_bank_rd_data_out_1_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22621 = _T_22620 | _T_22366; // @[Mux.scala 27:72]
  wire  _T_21606 = bht_rd_addr_hashed_f == 8'h3; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_3; // @[Reg.scala 27:20]
  wire [1:0] _T_22367 = _T_21606 ? bht_bank_rd_data_out_1_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22622 = _T_22621 | _T_22367; // @[Mux.scala 27:72]
  wire  _T_21609 = bht_rd_addr_hashed_f == 8'h4; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_4; // @[Reg.scala 27:20]
  wire [1:0] _T_22368 = _T_21609 ? bht_bank_rd_data_out_1_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22623 = _T_22622 | _T_22368; // @[Mux.scala 27:72]
  wire  _T_21612 = bht_rd_addr_hashed_f == 8'h5; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_5; // @[Reg.scala 27:20]
  wire [1:0] _T_22369 = _T_21612 ? bht_bank_rd_data_out_1_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22624 = _T_22623 | _T_22369; // @[Mux.scala 27:72]
  wire  _T_21615 = bht_rd_addr_hashed_f == 8'h6; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_6; // @[Reg.scala 27:20]
  wire [1:0] _T_22370 = _T_21615 ? bht_bank_rd_data_out_1_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22625 = _T_22624 | _T_22370; // @[Mux.scala 27:72]
  wire  _T_21618 = bht_rd_addr_hashed_f == 8'h7; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_7; // @[Reg.scala 27:20]
  wire [1:0] _T_22371 = _T_21618 ? bht_bank_rd_data_out_1_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22626 = _T_22625 | _T_22371; // @[Mux.scala 27:72]
  wire  _T_21621 = bht_rd_addr_hashed_f == 8'h8; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_8; // @[Reg.scala 27:20]
  wire [1:0] _T_22372 = _T_21621 ? bht_bank_rd_data_out_1_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22627 = _T_22626 | _T_22372; // @[Mux.scala 27:72]
  wire  _T_21624 = bht_rd_addr_hashed_f == 8'h9; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_9; // @[Reg.scala 27:20]
  wire [1:0] _T_22373 = _T_21624 ? bht_bank_rd_data_out_1_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22628 = _T_22627 | _T_22373; // @[Mux.scala 27:72]
  wire  _T_21627 = bht_rd_addr_hashed_f == 8'ha; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_10; // @[Reg.scala 27:20]
  wire [1:0] _T_22374 = _T_21627 ? bht_bank_rd_data_out_1_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22629 = _T_22628 | _T_22374; // @[Mux.scala 27:72]
  wire  _T_21630 = bht_rd_addr_hashed_f == 8'hb; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_11; // @[Reg.scala 27:20]
  wire [1:0] _T_22375 = _T_21630 ? bht_bank_rd_data_out_1_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22630 = _T_22629 | _T_22375; // @[Mux.scala 27:72]
  wire  _T_21633 = bht_rd_addr_hashed_f == 8'hc; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_12; // @[Reg.scala 27:20]
  wire [1:0] _T_22376 = _T_21633 ? bht_bank_rd_data_out_1_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22631 = _T_22630 | _T_22376; // @[Mux.scala 27:72]
  wire  _T_21636 = bht_rd_addr_hashed_f == 8'hd; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_13; // @[Reg.scala 27:20]
  wire [1:0] _T_22377 = _T_21636 ? bht_bank_rd_data_out_1_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22632 = _T_22631 | _T_22377; // @[Mux.scala 27:72]
  wire  _T_21639 = bht_rd_addr_hashed_f == 8'he; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_14; // @[Reg.scala 27:20]
  wire [1:0] _T_22378 = _T_21639 ? bht_bank_rd_data_out_1_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22633 = _T_22632 | _T_22378; // @[Mux.scala 27:72]
  wire  _T_21642 = bht_rd_addr_hashed_f == 8'hf; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_15; // @[Reg.scala 27:20]
  wire [1:0] _T_22379 = _T_21642 ? bht_bank_rd_data_out_1_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22634 = _T_22633 | _T_22379; // @[Mux.scala 27:72]
  wire  _T_21645 = bht_rd_addr_hashed_f == 8'h10; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_16; // @[Reg.scala 27:20]
  wire [1:0] _T_22380 = _T_21645 ? bht_bank_rd_data_out_1_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22635 = _T_22634 | _T_22380; // @[Mux.scala 27:72]
  wire  _T_21648 = bht_rd_addr_hashed_f == 8'h11; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_17; // @[Reg.scala 27:20]
  wire [1:0] _T_22381 = _T_21648 ? bht_bank_rd_data_out_1_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22636 = _T_22635 | _T_22381; // @[Mux.scala 27:72]
  wire  _T_21651 = bht_rd_addr_hashed_f == 8'h12; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_18; // @[Reg.scala 27:20]
  wire [1:0] _T_22382 = _T_21651 ? bht_bank_rd_data_out_1_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22637 = _T_22636 | _T_22382; // @[Mux.scala 27:72]
  wire  _T_21654 = bht_rd_addr_hashed_f == 8'h13; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_19; // @[Reg.scala 27:20]
  wire [1:0] _T_22383 = _T_21654 ? bht_bank_rd_data_out_1_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22638 = _T_22637 | _T_22383; // @[Mux.scala 27:72]
  wire  _T_21657 = bht_rd_addr_hashed_f == 8'h14; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_20; // @[Reg.scala 27:20]
  wire [1:0] _T_22384 = _T_21657 ? bht_bank_rd_data_out_1_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22639 = _T_22638 | _T_22384; // @[Mux.scala 27:72]
  wire  _T_21660 = bht_rd_addr_hashed_f == 8'h15; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_21; // @[Reg.scala 27:20]
  wire [1:0] _T_22385 = _T_21660 ? bht_bank_rd_data_out_1_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22640 = _T_22639 | _T_22385; // @[Mux.scala 27:72]
  wire  _T_21663 = bht_rd_addr_hashed_f == 8'h16; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_22; // @[Reg.scala 27:20]
  wire [1:0] _T_22386 = _T_21663 ? bht_bank_rd_data_out_1_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22641 = _T_22640 | _T_22386; // @[Mux.scala 27:72]
  wire  _T_21666 = bht_rd_addr_hashed_f == 8'h17; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_23; // @[Reg.scala 27:20]
  wire [1:0] _T_22387 = _T_21666 ? bht_bank_rd_data_out_1_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22642 = _T_22641 | _T_22387; // @[Mux.scala 27:72]
  wire  _T_21669 = bht_rd_addr_hashed_f == 8'h18; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_24; // @[Reg.scala 27:20]
  wire [1:0] _T_22388 = _T_21669 ? bht_bank_rd_data_out_1_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22643 = _T_22642 | _T_22388; // @[Mux.scala 27:72]
  wire  _T_21672 = bht_rd_addr_hashed_f == 8'h19; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_25; // @[Reg.scala 27:20]
  wire [1:0] _T_22389 = _T_21672 ? bht_bank_rd_data_out_1_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22644 = _T_22643 | _T_22389; // @[Mux.scala 27:72]
  wire  _T_21675 = bht_rd_addr_hashed_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_26; // @[Reg.scala 27:20]
  wire [1:0] _T_22390 = _T_21675 ? bht_bank_rd_data_out_1_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22645 = _T_22644 | _T_22390; // @[Mux.scala 27:72]
  wire  _T_21678 = bht_rd_addr_hashed_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_27; // @[Reg.scala 27:20]
  wire [1:0] _T_22391 = _T_21678 ? bht_bank_rd_data_out_1_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22646 = _T_22645 | _T_22391; // @[Mux.scala 27:72]
  wire  _T_21681 = bht_rd_addr_hashed_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_28; // @[Reg.scala 27:20]
  wire [1:0] _T_22392 = _T_21681 ? bht_bank_rd_data_out_1_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22647 = _T_22646 | _T_22392; // @[Mux.scala 27:72]
  wire  _T_21684 = bht_rd_addr_hashed_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_29; // @[Reg.scala 27:20]
  wire [1:0] _T_22393 = _T_21684 ? bht_bank_rd_data_out_1_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22648 = _T_22647 | _T_22393; // @[Mux.scala 27:72]
  wire  _T_21687 = bht_rd_addr_hashed_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_30; // @[Reg.scala 27:20]
  wire [1:0] _T_22394 = _T_21687 ? bht_bank_rd_data_out_1_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22649 = _T_22648 | _T_22394; // @[Mux.scala 27:72]
  wire  _T_21690 = bht_rd_addr_hashed_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_31; // @[Reg.scala 27:20]
  wire [1:0] _T_22395 = _T_21690 ? bht_bank_rd_data_out_1_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22650 = _T_22649 | _T_22395; // @[Mux.scala 27:72]
  wire  _T_21693 = bht_rd_addr_hashed_f == 8'h20; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_32; // @[Reg.scala 27:20]
  wire [1:0] _T_22396 = _T_21693 ? bht_bank_rd_data_out_1_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22651 = _T_22650 | _T_22396; // @[Mux.scala 27:72]
  wire  _T_21696 = bht_rd_addr_hashed_f == 8'h21; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_33; // @[Reg.scala 27:20]
  wire [1:0] _T_22397 = _T_21696 ? bht_bank_rd_data_out_1_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22652 = _T_22651 | _T_22397; // @[Mux.scala 27:72]
  wire  _T_21699 = bht_rd_addr_hashed_f == 8'h22; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_34; // @[Reg.scala 27:20]
  wire [1:0] _T_22398 = _T_21699 ? bht_bank_rd_data_out_1_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22653 = _T_22652 | _T_22398; // @[Mux.scala 27:72]
  wire  _T_21702 = bht_rd_addr_hashed_f == 8'h23; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_35; // @[Reg.scala 27:20]
  wire [1:0] _T_22399 = _T_21702 ? bht_bank_rd_data_out_1_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22654 = _T_22653 | _T_22399; // @[Mux.scala 27:72]
  wire  _T_21705 = bht_rd_addr_hashed_f == 8'h24; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_36; // @[Reg.scala 27:20]
  wire [1:0] _T_22400 = _T_21705 ? bht_bank_rd_data_out_1_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22655 = _T_22654 | _T_22400; // @[Mux.scala 27:72]
  wire  _T_21708 = bht_rd_addr_hashed_f == 8'h25; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_37; // @[Reg.scala 27:20]
  wire [1:0] _T_22401 = _T_21708 ? bht_bank_rd_data_out_1_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22656 = _T_22655 | _T_22401; // @[Mux.scala 27:72]
  wire  _T_21711 = bht_rd_addr_hashed_f == 8'h26; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_38; // @[Reg.scala 27:20]
  wire [1:0] _T_22402 = _T_21711 ? bht_bank_rd_data_out_1_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22657 = _T_22656 | _T_22402; // @[Mux.scala 27:72]
  wire  _T_21714 = bht_rd_addr_hashed_f == 8'h27; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_39; // @[Reg.scala 27:20]
  wire [1:0] _T_22403 = _T_21714 ? bht_bank_rd_data_out_1_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22658 = _T_22657 | _T_22403; // @[Mux.scala 27:72]
  wire  _T_21717 = bht_rd_addr_hashed_f == 8'h28; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_40; // @[Reg.scala 27:20]
  wire [1:0] _T_22404 = _T_21717 ? bht_bank_rd_data_out_1_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22659 = _T_22658 | _T_22404; // @[Mux.scala 27:72]
  wire  _T_21720 = bht_rd_addr_hashed_f == 8'h29; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_41; // @[Reg.scala 27:20]
  wire [1:0] _T_22405 = _T_21720 ? bht_bank_rd_data_out_1_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22660 = _T_22659 | _T_22405; // @[Mux.scala 27:72]
  wire  _T_21723 = bht_rd_addr_hashed_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_42; // @[Reg.scala 27:20]
  wire [1:0] _T_22406 = _T_21723 ? bht_bank_rd_data_out_1_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22661 = _T_22660 | _T_22406; // @[Mux.scala 27:72]
  wire  _T_21726 = bht_rd_addr_hashed_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_43; // @[Reg.scala 27:20]
  wire [1:0] _T_22407 = _T_21726 ? bht_bank_rd_data_out_1_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22662 = _T_22661 | _T_22407; // @[Mux.scala 27:72]
  wire  _T_21729 = bht_rd_addr_hashed_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_44; // @[Reg.scala 27:20]
  wire [1:0] _T_22408 = _T_21729 ? bht_bank_rd_data_out_1_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22663 = _T_22662 | _T_22408; // @[Mux.scala 27:72]
  wire  _T_21732 = bht_rd_addr_hashed_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_45; // @[Reg.scala 27:20]
  wire [1:0] _T_22409 = _T_21732 ? bht_bank_rd_data_out_1_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22664 = _T_22663 | _T_22409; // @[Mux.scala 27:72]
  wire  _T_21735 = bht_rd_addr_hashed_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_46; // @[Reg.scala 27:20]
  wire [1:0] _T_22410 = _T_21735 ? bht_bank_rd_data_out_1_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22665 = _T_22664 | _T_22410; // @[Mux.scala 27:72]
  wire  _T_21738 = bht_rd_addr_hashed_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_47; // @[Reg.scala 27:20]
  wire [1:0] _T_22411 = _T_21738 ? bht_bank_rd_data_out_1_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22666 = _T_22665 | _T_22411; // @[Mux.scala 27:72]
  wire  _T_21741 = bht_rd_addr_hashed_f == 8'h30; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_48; // @[Reg.scala 27:20]
  wire [1:0] _T_22412 = _T_21741 ? bht_bank_rd_data_out_1_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22667 = _T_22666 | _T_22412; // @[Mux.scala 27:72]
  wire  _T_21744 = bht_rd_addr_hashed_f == 8'h31; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_49; // @[Reg.scala 27:20]
  wire [1:0] _T_22413 = _T_21744 ? bht_bank_rd_data_out_1_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22668 = _T_22667 | _T_22413; // @[Mux.scala 27:72]
  wire  _T_21747 = bht_rd_addr_hashed_f == 8'h32; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_50; // @[Reg.scala 27:20]
  wire [1:0] _T_22414 = _T_21747 ? bht_bank_rd_data_out_1_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22669 = _T_22668 | _T_22414; // @[Mux.scala 27:72]
  wire  _T_21750 = bht_rd_addr_hashed_f == 8'h33; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_51; // @[Reg.scala 27:20]
  wire [1:0] _T_22415 = _T_21750 ? bht_bank_rd_data_out_1_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22670 = _T_22669 | _T_22415; // @[Mux.scala 27:72]
  wire  _T_21753 = bht_rd_addr_hashed_f == 8'h34; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_52; // @[Reg.scala 27:20]
  wire [1:0] _T_22416 = _T_21753 ? bht_bank_rd_data_out_1_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22671 = _T_22670 | _T_22416; // @[Mux.scala 27:72]
  wire  _T_21756 = bht_rd_addr_hashed_f == 8'h35; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_53; // @[Reg.scala 27:20]
  wire [1:0] _T_22417 = _T_21756 ? bht_bank_rd_data_out_1_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22672 = _T_22671 | _T_22417; // @[Mux.scala 27:72]
  wire  _T_21759 = bht_rd_addr_hashed_f == 8'h36; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_54; // @[Reg.scala 27:20]
  wire [1:0] _T_22418 = _T_21759 ? bht_bank_rd_data_out_1_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22673 = _T_22672 | _T_22418; // @[Mux.scala 27:72]
  wire  _T_21762 = bht_rd_addr_hashed_f == 8'h37; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_55; // @[Reg.scala 27:20]
  wire [1:0] _T_22419 = _T_21762 ? bht_bank_rd_data_out_1_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22674 = _T_22673 | _T_22419; // @[Mux.scala 27:72]
  wire  _T_21765 = bht_rd_addr_hashed_f == 8'h38; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_56; // @[Reg.scala 27:20]
  wire [1:0] _T_22420 = _T_21765 ? bht_bank_rd_data_out_1_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22675 = _T_22674 | _T_22420; // @[Mux.scala 27:72]
  wire  _T_21768 = bht_rd_addr_hashed_f == 8'h39; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_57; // @[Reg.scala 27:20]
  wire [1:0] _T_22421 = _T_21768 ? bht_bank_rd_data_out_1_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22676 = _T_22675 | _T_22421; // @[Mux.scala 27:72]
  wire  _T_21771 = bht_rd_addr_hashed_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_58; // @[Reg.scala 27:20]
  wire [1:0] _T_22422 = _T_21771 ? bht_bank_rd_data_out_1_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22677 = _T_22676 | _T_22422; // @[Mux.scala 27:72]
  wire  _T_21774 = bht_rd_addr_hashed_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_59; // @[Reg.scala 27:20]
  wire [1:0] _T_22423 = _T_21774 ? bht_bank_rd_data_out_1_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22678 = _T_22677 | _T_22423; // @[Mux.scala 27:72]
  wire  _T_21777 = bht_rd_addr_hashed_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_60; // @[Reg.scala 27:20]
  wire [1:0] _T_22424 = _T_21777 ? bht_bank_rd_data_out_1_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22679 = _T_22678 | _T_22424; // @[Mux.scala 27:72]
  wire  _T_21780 = bht_rd_addr_hashed_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_61; // @[Reg.scala 27:20]
  wire [1:0] _T_22425 = _T_21780 ? bht_bank_rd_data_out_1_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22680 = _T_22679 | _T_22425; // @[Mux.scala 27:72]
  wire  _T_21783 = bht_rd_addr_hashed_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_62; // @[Reg.scala 27:20]
  wire [1:0] _T_22426 = _T_21783 ? bht_bank_rd_data_out_1_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22681 = _T_22680 | _T_22426; // @[Mux.scala 27:72]
  wire  _T_21786 = bht_rd_addr_hashed_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_63; // @[Reg.scala 27:20]
  wire [1:0] _T_22427 = _T_21786 ? bht_bank_rd_data_out_1_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22682 = _T_22681 | _T_22427; // @[Mux.scala 27:72]
  wire  _T_21789 = bht_rd_addr_hashed_f == 8'h40; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_64; // @[Reg.scala 27:20]
  wire [1:0] _T_22428 = _T_21789 ? bht_bank_rd_data_out_1_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22683 = _T_22682 | _T_22428; // @[Mux.scala 27:72]
  wire  _T_21792 = bht_rd_addr_hashed_f == 8'h41; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_65; // @[Reg.scala 27:20]
  wire [1:0] _T_22429 = _T_21792 ? bht_bank_rd_data_out_1_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22684 = _T_22683 | _T_22429; // @[Mux.scala 27:72]
  wire  _T_21795 = bht_rd_addr_hashed_f == 8'h42; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_66; // @[Reg.scala 27:20]
  wire [1:0] _T_22430 = _T_21795 ? bht_bank_rd_data_out_1_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22685 = _T_22684 | _T_22430; // @[Mux.scala 27:72]
  wire  _T_21798 = bht_rd_addr_hashed_f == 8'h43; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_67; // @[Reg.scala 27:20]
  wire [1:0] _T_22431 = _T_21798 ? bht_bank_rd_data_out_1_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22686 = _T_22685 | _T_22431; // @[Mux.scala 27:72]
  wire  _T_21801 = bht_rd_addr_hashed_f == 8'h44; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_68; // @[Reg.scala 27:20]
  wire [1:0] _T_22432 = _T_21801 ? bht_bank_rd_data_out_1_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22687 = _T_22686 | _T_22432; // @[Mux.scala 27:72]
  wire  _T_21804 = bht_rd_addr_hashed_f == 8'h45; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_69; // @[Reg.scala 27:20]
  wire [1:0] _T_22433 = _T_21804 ? bht_bank_rd_data_out_1_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22688 = _T_22687 | _T_22433; // @[Mux.scala 27:72]
  wire  _T_21807 = bht_rd_addr_hashed_f == 8'h46; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_70; // @[Reg.scala 27:20]
  wire [1:0] _T_22434 = _T_21807 ? bht_bank_rd_data_out_1_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22689 = _T_22688 | _T_22434; // @[Mux.scala 27:72]
  wire  _T_21810 = bht_rd_addr_hashed_f == 8'h47; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_71; // @[Reg.scala 27:20]
  wire [1:0] _T_22435 = _T_21810 ? bht_bank_rd_data_out_1_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22690 = _T_22689 | _T_22435; // @[Mux.scala 27:72]
  wire  _T_21813 = bht_rd_addr_hashed_f == 8'h48; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_72; // @[Reg.scala 27:20]
  wire [1:0] _T_22436 = _T_21813 ? bht_bank_rd_data_out_1_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22691 = _T_22690 | _T_22436; // @[Mux.scala 27:72]
  wire  _T_21816 = bht_rd_addr_hashed_f == 8'h49; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_73; // @[Reg.scala 27:20]
  wire [1:0] _T_22437 = _T_21816 ? bht_bank_rd_data_out_1_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22692 = _T_22691 | _T_22437; // @[Mux.scala 27:72]
  wire  _T_21819 = bht_rd_addr_hashed_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_74; // @[Reg.scala 27:20]
  wire [1:0] _T_22438 = _T_21819 ? bht_bank_rd_data_out_1_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22693 = _T_22692 | _T_22438; // @[Mux.scala 27:72]
  wire  _T_21822 = bht_rd_addr_hashed_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_75; // @[Reg.scala 27:20]
  wire [1:0] _T_22439 = _T_21822 ? bht_bank_rd_data_out_1_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22694 = _T_22693 | _T_22439; // @[Mux.scala 27:72]
  wire  _T_21825 = bht_rd_addr_hashed_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_76; // @[Reg.scala 27:20]
  wire [1:0] _T_22440 = _T_21825 ? bht_bank_rd_data_out_1_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22695 = _T_22694 | _T_22440; // @[Mux.scala 27:72]
  wire  _T_21828 = bht_rd_addr_hashed_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_77; // @[Reg.scala 27:20]
  wire [1:0] _T_22441 = _T_21828 ? bht_bank_rd_data_out_1_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22696 = _T_22695 | _T_22441; // @[Mux.scala 27:72]
  wire  _T_21831 = bht_rd_addr_hashed_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_78; // @[Reg.scala 27:20]
  wire [1:0] _T_22442 = _T_21831 ? bht_bank_rd_data_out_1_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22697 = _T_22696 | _T_22442; // @[Mux.scala 27:72]
  wire  _T_21834 = bht_rd_addr_hashed_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_79; // @[Reg.scala 27:20]
  wire [1:0] _T_22443 = _T_21834 ? bht_bank_rd_data_out_1_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22698 = _T_22697 | _T_22443; // @[Mux.scala 27:72]
  wire  _T_21837 = bht_rd_addr_hashed_f == 8'h50; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_80; // @[Reg.scala 27:20]
  wire [1:0] _T_22444 = _T_21837 ? bht_bank_rd_data_out_1_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22699 = _T_22698 | _T_22444; // @[Mux.scala 27:72]
  wire  _T_21840 = bht_rd_addr_hashed_f == 8'h51; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_81; // @[Reg.scala 27:20]
  wire [1:0] _T_22445 = _T_21840 ? bht_bank_rd_data_out_1_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22700 = _T_22699 | _T_22445; // @[Mux.scala 27:72]
  wire  _T_21843 = bht_rd_addr_hashed_f == 8'h52; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_82; // @[Reg.scala 27:20]
  wire [1:0] _T_22446 = _T_21843 ? bht_bank_rd_data_out_1_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22701 = _T_22700 | _T_22446; // @[Mux.scala 27:72]
  wire  _T_21846 = bht_rd_addr_hashed_f == 8'h53; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_83; // @[Reg.scala 27:20]
  wire [1:0] _T_22447 = _T_21846 ? bht_bank_rd_data_out_1_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22702 = _T_22701 | _T_22447; // @[Mux.scala 27:72]
  wire  _T_21849 = bht_rd_addr_hashed_f == 8'h54; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_84; // @[Reg.scala 27:20]
  wire [1:0] _T_22448 = _T_21849 ? bht_bank_rd_data_out_1_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22703 = _T_22702 | _T_22448; // @[Mux.scala 27:72]
  wire  _T_21852 = bht_rd_addr_hashed_f == 8'h55; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_85; // @[Reg.scala 27:20]
  wire [1:0] _T_22449 = _T_21852 ? bht_bank_rd_data_out_1_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22704 = _T_22703 | _T_22449; // @[Mux.scala 27:72]
  wire  _T_21855 = bht_rd_addr_hashed_f == 8'h56; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_86; // @[Reg.scala 27:20]
  wire [1:0] _T_22450 = _T_21855 ? bht_bank_rd_data_out_1_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22705 = _T_22704 | _T_22450; // @[Mux.scala 27:72]
  wire  _T_21858 = bht_rd_addr_hashed_f == 8'h57; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_87; // @[Reg.scala 27:20]
  wire [1:0] _T_22451 = _T_21858 ? bht_bank_rd_data_out_1_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22706 = _T_22705 | _T_22451; // @[Mux.scala 27:72]
  wire  _T_21861 = bht_rd_addr_hashed_f == 8'h58; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_88; // @[Reg.scala 27:20]
  wire [1:0] _T_22452 = _T_21861 ? bht_bank_rd_data_out_1_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22707 = _T_22706 | _T_22452; // @[Mux.scala 27:72]
  wire  _T_21864 = bht_rd_addr_hashed_f == 8'h59; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_89; // @[Reg.scala 27:20]
  wire [1:0] _T_22453 = _T_21864 ? bht_bank_rd_data_out_1_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22708 = _T_22707 | _T_22453; // @[Mux.scala 27:72]
  wire  _T_21867 = bht_rd_addr_hashed_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_90; // @[Reg.scala 27:20]
  wire [1:0] _T_22454 = _T_21867 ? bht_bank_rd_data_out_1_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22709 = _T_22708 | _T_22454; // @[Mux.scala 27:72]
  wire  _T_21870 = bht_rd_addr_hashed_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_91; // @[Reg.scala 27:20]
  wire [1:0] _T_22455 = _T_21870 ? bht_bank_rd_data_out_1_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22710 = _T_22709 | _T_22455; // @[Mux.scala 27:72]
  wire  _T_21873 = bht_rd_addr_hashed_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_92; // @[Reg.scala 27:20]
  wire [1:0] _T_22456 = _T_21873 ? bht_bank_rd_data_out_1_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22711 = _T_22710 | _T_22456; // @[Mux.scala 27:72]
  wire  _T_21876 = bht_rd_addr_hashed_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_93; // @[Reg.scala 27:20]
  wire [1:0] _T_22457 = _T_21876 ? bht_bank_rd_data_out_1_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22712 = _T_22711 | _T_22457; // @[Mux.scala 27:72]
  wire  _T_21879 = bht_rd_addr_hashed_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_94; // @[Reg.scala 27:20]
  wire [1:0] _T_22458 = _T_21879 ? bht_bank_rd_data_out_1_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22713 = _T_22712 | _T_22458; // @[Mux.scala 27:72]
  wire  _T_21882 = bht_rd_addr_hashed_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_95; // @[Reg.scala 27:20]
  wire [1:0] _T_22459 = _T_21882 ? bht_bank_rd_data_out_1_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22714 = _T_22713 | _T_22459; // @[Mux.scala 27:72]
  wire  _T_21885 = bht_rd_addr_hashed_f == 8'h60; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_96; // @[Reg.scala 27:20]
  wire [1:0] _T_22460 = _T_21885 ? bht_bank_rd_data_out_1_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22715 = _T_22714 | _T_22460; // @[Mux.scala 27:72]
  wire  _T_21888 = bht_rd_addr_hashed_f == 8'h61; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_97; // @[Reg.scala 27:20]
  wire [1:0] _T_22461 = _T_21888 ? bht_bank_rd_data_out_1_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22716 = _T_22715 | _T_22461; // @[Mux.scala 27:72]
  wire  _T_21891 = bht_rd_addr_hashed_f == 8'h62; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_98; // @[Reg.scala 27:20]
  wire [1:0] _T_22462 = _T_21891 ? bht_bank_rd_data_out_1_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22717 = _T_22716 | _T_22462; // @[Mux.scala 27:72]
  wire  _T_21894 = bht_rd_addr_hashed_f == 8'h63; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_99; // @[Reg.scala 27:20]
  wire [1:0] _T_22463 = _T_21894 ? bht_bank_rd_data_out_1_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22718 = _T_22717 | _T_22463; // @[Mux.scala 27:72]
  wire  _T_21897 = bht_rd_addr_hashed_f == 8'h64; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_100; // @[Reg.scala 27:20]
  wire [1:0] _T_22464 = _T_21897 ? bht_bank_rd_data_out_1_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22719 = _T_22718 | _T_22464; // @[Mux.scala 27:72]
  wire  _T_21900 = bht_rd_addr_hashed_f == 8'h65; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_101; // @[Reg.scala 27:20]
  wire [1:0] _T_22465 = _T_21900 ? bht_bank_rd_data_out_1_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22720 = _T_22719 | _T_22465; // @[Mux.scala 27:72]
  wire  _T_21903 = bht_rd_addr_hashed_f == 8'h66; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_102; // @[Reg.scala 27:20]
  wire [1:0] _T_22466 = _T_21903 ? bht_bank_rd_data_out_1_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22721 = _T_22720 | _T_22466; // @[Mux.scala 27:72]
  wire  _T_21906 = bht_rd_addr_hashed_f == 8'h67; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_103; // @[Reg.scala 27:20]
  wire [1:0] _T_22467 = _T_21906 ? bht_bank_rd_data_out_1_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22722 = _T_22721 | _T_22467; // @[Mux.scala 27:72]
  wire  _T_21909 = bht_rd_addr_hashed_f == 8'h68; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_104; // @[Reg.scala 27:20]
  wire [1:0] _T_22468 = _T_21909 ? bht_bank_rd_data_out_1_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22723 = _T_22722 | _T_22468; // @[Mux.scala 27:72]
  wire  _T_21912 = bht_rd_addr_hashed_f == 8'h69; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_105; // @[Reg.scala 27:20]
  wire [1:0] _T_22469 = _T_21912 ? bht_bank_rd_data_out_1_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22724 = _T_22723 | _T_22469; // @[Mux.scala 27:72]
  wire  _T_21915 = bht_rd_addr_hashed_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_106; // @[Reg.scala 27:20]
  wire [1:0] _T_22470 = _T_21915 ? bht_bank_rd_data_out_1_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22725 = _T_22724 | _T_22470; // @[Mux.scala 27:72]
  wire  _T_21918 = bht_rd_addr_hashed_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_107; // @[Reg.scala 27:20]
  wire [1:0] _T_22471 = _T_21918 ? bht_bank_rd_data_out_1_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22726 = _T_22725 | _T_22471; // @[Mux.scala 27:72]
  wire  _T_21921 = bht_rd_addr_hashed_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_108; // @[Reg.scala 27:20]
  wire [1:0] _T_22472 = _T_21921 ? bht_bank_rd_data_out_1_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22727 = _T_22726 | _T_22472; // @[Mux.scala 27:72]
  wire  _T_21924 = bht_rd_addr_hashed_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_109; // @[Reg.scala 27:20]
  wire [1:0] _T_22473 = _T_21924 ? bht_bank_rd_data_out_1_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22728 = _T_22727 | _T_22473; // @[Mux.scala 27:72]
  wire  _T_21927 = bht_rd_addr_hashed_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_110; // @[Reg.scala 27:20]
  wire [1:0] _T_22474 = _T_21927 ? bht_bank_rd_data_out_1_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22729 = _T_22728 | _T_22474; // @[Mux.scala 27:72]
  wire  _T_21930 = bht_rd_addr_hashed_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_111; // @[Reg.scala 27:20]
  wire [1:0] _T_22475 = _T_21930 ? bht_bank_rd_data_out_1_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22730 = _T_22729 | _T_22475; // @[Mux.scala 27:72]
  wire  _T_21933 = bht_rd_addr_hashed_f == 8'h70; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_112; // @[Reg.scala 27:20]
  wire [1:0] _T_22476 = _T_21933 ? bht_bank_rd_data_out_1_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22731 = _T_22730 | _T_22476; // @[Mux.scala 27:72]
  wire  _T_21936 = bht_rd_addr_hashed_f == 8'h71; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_113; // @[Reg.scala 27:20]
  wire [1:0] _T_22477 = _T_21936 ? bht_bank_rd_data_out_1_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22732 = _T_22731 | _T_22477; // @[Mux.scala 27:72]
  wire  _T_21939 = bht_rd_addr_hashed_f == 8'h72; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_114; // @[Reg.scala 27:20]
  wire [1:0] _T_22478 = _T_21939 ? bht_bank_rd_data_out_1_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22733 = _T_22732 | _T_22478; // @[Mux.scala 27:72]
  wire  _T_21942 = bht_rd_addr_hashed_f == 8'h73; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_115; // @[Reg.scala 27:20]
  wire [1:0] _T_22479 = _T_21942 ? bht_bank_rd_data_out_1_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22734 = _T_22733 | _T_22479; // @[Mux.scala 27:72]
  wire  _T_21945 = bht_rd_addr_hashed_f == 8'h74; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_116; // @[Reg.scala 27:20]
  wire [1:0] _T_22480 = _T_21945 ? bht_bank_rd_data_out_1_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22735 = _T_22734 | _T_22480; // @[Mux.scala 27:72]
  wire  _T_21948 = bht_rd_addr_hashed_f == 8'h75; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_117; // @[Reg.scala 27:20]
  wire [1:0] _T_22481 = _T_21948 ? bht_bank_rd_data_out_1_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22736 = _T_22735 | _T_22481; // @[Mux.scala 27:72]
  wire  _T_21951 = bht_rd_addr_hashed_f == 8'h76; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_118; // @[Reg.scala 27:20]
  wire [1:0] _T_22482 = _T_21951 ? bht_bank_rd_data_out_1_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22737 = _T_22736 | _T_22482; // @[Mux.scala 27:72]
  wire  _T_21954 = bht_rd_addr_hashed_f == 8'h77; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_119; // @[Reg.scala 27:20]
  wire [1:0] _T_22483 = _T_21954 ? bht_bank_rd_data_out_1_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22738 = _T_22737 | _T_22483; // @[Mux.scala 27:72]
  wire  _T_21957 = bht_rd_addr_hashed_f == 8'h78; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_120; // @[Reg.scala 27:20]
  wire [1:0] _T_22484 = _T_21957 ? bht_bank_rd_data_out_1_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22739 = _T_22738 | _T_22484; // @[Mux.scala 27:72]
  wire  _T_21960 = bht_rd_addr_hashed_f == 8'h79; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_121; // @[Reg.scala 27:20]
  wire [1:0] _T_22485 = _T_21960 ? bht_bank_rd_data_out_1_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22740 = _T_22739 | _T_22485; // @[Mux.scala 27:72]
  wire  _T_21963 = bht_rd_addr_hashed_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_122; // @[Reg.scala 27:20]
  wire [1:0] _T_22486 = _T_21963 ? bht_bank_rd_data_out_1_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22741 = _T_22740 | _T_22486; // @[Mux.scala 27:72]
  wire  _T_21966 = bht_rd_addr_hashed_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_123; // @[Reg.scala 27:20]
  wire [1:0] _T_22487 = _T_21966 ? bht_bank_rd_data_out_1_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22742 = _T_22741 | _T_22487; // @[Mux.scala 27:72]
  wire  _T_21969 = bht_rd_addr_hashed_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_124; // @[Reg.scala 27:20]
  wire [1:0] _T_22488 = _T_21969 ? bht_bank_rd_data_out_1_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22743 = _T_22742 | _T_22488; // @[Mux.scala 27:72]
  wire  _T_21972 = bht_rd_addr_hashed_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_125; // @[Reg.scala 27:20]
  wire [1:0] _T_22489 = _T_21972 ? bht_bank_rd_data_out_1_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22744 = _T_22743 | _T_22489; // @[Mux.scala 27:72]
  wire  _T_21975 = bht_rd_addr_hashed_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_126; // @[Reg.scala 27:20]
  wire [1:0] _T_22490 = _T_21975 ? bht_bank_rd_data_out_1_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22745 = _T_22744 | _T_22490; // @[Mux.scala 27:72]
  wire  _T_21978 = bht_rd_addr_hashed_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_127; // @[Reg.scala 27:20]
  wire [1:0] _T_22491 = _T_21978 ? bht_bank_rd_data_out_1_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22746 = _T_22745 | _T_22491; // @[Mux.scala 27:72]
  wire  _T_21981 = bht_rd_addr_hashed_f == 8'h80; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_128; // @[Reg.scala 27:20]
  wire [1:0] _T_22492 = _T_21981 ? bht_bank_rd_data_out_1_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22747 = _T_22746 | _T_22492; // @[Mux.scala 27:72]
  wire  _T_21984 = bht_rd_addr_hashed_f == 8'h81; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_129; // @[Reg.scala 27:20]
  wire [1:0] _T_22493 = _T_21984 ? bht_bank_rd_data_out_1_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22748 = _T_22747 | _T_22493; // @[Mux.scala 27:72]
  wire  _T_21987 = bht_rd_addr_hashed_f == 8'h82; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_130; // @[Reg.scala 27:20]
  wire [1:0] _T_22494 = _T_21987 ? bht_bank_rd_data_out_1_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22749 = _T_22748 | _T_22494; // @[Mux.scala 27:72]
  wire  _T_21990 = bht_rd_addr_hashed_f == 8'h83; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_131; // @[Reg.scala 27:20]
  wire [1:0] _T_22495 = _T_21990 ? bht_bank_rd_data_out_1_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22750 = _T_22749 | _T_22495; // @[Mux.scala 27:72]
  wire  _T_21993 = bht_rd_addr_hashed_f == 8'h84; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_132; // @[Reg.scala 27:20]
  wire [1:0] _T_22496 = _T_21993 ? bht_bank_rd_data_out_1_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22751 = _T_22750 | _T_22496; // @[Mux.scala 27:72]
  wire  _T_21996 = bht_rd_addr_hashed_f == 8'h85; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_133; // @[Reg.scala 27:20]
  wire [1:0] _T_22497 = _T_21996 ? bht_bank_rd_data_out_1_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22752 = _T_22751 | _T_22497; // @[Mux.scala 27:72]
  wire  _T_21999 = bht_rd_addr_hashed_f == 8'h86; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_134; // @[Reg.scala 27:20]
  wire [1:0] _T_22498 = _T_21999 ? bht_bank_rd_data_out_1_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22753 = _T_22752 | _T_22498; // @[Mux.scala 27:72]
  wire  _T_22002 = bht_rd_addr_hashed_f == 8'h87; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_135; // @[Reg.scala 27:20]
  wire [1:0] _T_22499 = _T_22002 ? bht_bank_rd_data_out_1_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22754 = _T_22753 | _T_22499; // @[Mux.scala 27:72]
  wire  _T_22005 = bht_rd_addr_hashed_f == 8'h88; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_136; // @[Reg.scala 27:20]
  wire [1:0] _T_22500 = _T_22005 ? bht_bank_rd_data_out_1_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22755 = _T_22754 | _T_22500; // @[Mux.scala 27:72]
  wire  _T_22008 = bht_rd_addr_hashed_f == 8'h89; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_137; // @[Reg.scala 27:20]
  wire [1:0] _T_22501 = _T_22008 ? bht_bank_rd_data_out_1_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22756 = _T_22755 | _T_22501; // @[Mux.scala 27:72]
  wire  _T_22011 = bht_rd_addr_hashed_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_138; // @[Reg.scala 27:20]
  wire [1:0] _T_22502 = _T_22011 ? bht_bank_rd_data_out_1_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22757 = _T_22756 | _T_22502; // @[Mux.scala 27:72]
  wire  _T_22014 = bht_rd_addr_hashed_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_139; // @[Reg.scala 27:20]
  wire [1:0] _T_22503 = _T_22014 ? bht_bank_rd_data_out_1_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22758 = _T_22757 | _T_22503; // @[Mux.scala 27:72]
  wire  _T_22017 = bht_rd_addr_hashed_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_140; // @[Reg.scala 27:20]
  wire [1:0] _T_22504 = _T_22017 ? bht_bank_rd_data_out_1_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22759 = _T_22758 | _T_22504; // @[Mux.scala 27:72]
  wire  _T_22020 = bht_rd_addr_hashed_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_141; // @[Reg.scala 27:20]
  wire [1:0] _T_22505 = _T_22020 ? bht_bank_rd_data_out_1_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22760 = _T_22759 | _T_22505; // @[Mux.scala 27:72]
  wire  _T_22023 = bht_rd_addr_hashed_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_142; // @[Reg.scala 27:20]
  wire [1:0] _T_22506 = _T_22023 ? bht_bank_rd_data_out_1_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22761 = _T_22760 | _T_22506; // @[Mux.scala 27:72]
  wire  _T_22026 = bht_rd_addr_hashed_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_143; // @[Reg.scala 27:20]
  wire [1:0] _T_22507 = _T_22026 ? bht_bank_rd_data_out_1_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22762 = _T_22761 | _T_22507; // @[Mux.scala 27:72]
  wire  _T_22029 = bht_rd_addr_hashed_f == 8'h90; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_144; // @[Reg.scala 27:20]
  wire [1:0] _T_22508 = _T_22029 ? bht_bank_rd_data_out_1_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22763 = _T_22762 | _T_22508; // @[Mux.scala 27:72]
  wire  _T_22032 = bht_rd_addr_hashed_f == 8'h91; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_145; // @[Reg.scala 27:20]
  wire [1:0] _T_22509 = _T_22032 ? bht_bank_rd_data_out_1_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22764 = _T_22763 | _T_22509; // @[Mux.scala 27:72]
  wire  _T_22035 = bht_rd_addr_hashed_f == 8'h92; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_146; // @[Reg.scala 27:20]
  wire [1:0] _T_22510 = _T_22035 ? bht_bank_rd_data_out_1_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22765 = _T_22764 | _T_22510; // @[Mux.scala 27:72]
  wire  _T_22038 = bht_rd_addr_hashed_f == 8'h93; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_147; // @[Reg.scala 27:20]
  wire [1:0] _T_22511 = _T_22038 ? bht_bank_rd_data_out_1_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22766 = _T_22765 | _T_22511; // @[Mux.scala 27:72]
  wire  _T_22041 = bht_rd_addr_hashed_f == 8'h94; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_148; // @[Reg.scala 27:20]
  wire [1:0] _T_22512 = _T_22041 ? bht_bank_rd_data_out_1_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22767 = _T_22766 | _T_22512; // @[Mux.scala 27:72]
  wire  _T_22044 = bht_rd_addr_hashed_f == 8'h95; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_149; // @[Reg.scala 27:20]
  wire [1:0] _T_22513 = _T_22044 ? bht_bank_rd_data_out_1_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22768 = _T_22767 | _T_22513; // @[Mux.scala 27:72]
  wire  _T_22047 = bht_rd_addr_hashed_f == 8'h96; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_150; // @[Reg.scala 27:20]
  wire [1:0] _T_22514 = _T_22047 ? bht_bank_rd_data_out_1_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22769 = _T_22768 | _T_22514; // @[Mux.scala 27:72]
  wire  _T_22050 = bht_rd_addr_hashed_f == 8'h97; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_151; // @[Reg.scala 27:20]
  wire [1:0] _T_22515 = _T_22050 ? bht_bank_rd_data_out_1_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22770 = _T_22769 | _T_22515; // @[Mux.scala 27:72]
  wire  _T_22053 = bht_rd_addr_hashed_f == 8'h98; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_152; // @[Reg.scala 27:20]
  wire [1:0] _T_22516 = _T_22053 ? bht_bank_rd_data_out_1_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22771 = _T_22770 | _T_22516; // @[Mux.scala 27:72]
  wire  _T_22056 = bht_rd_addr_hashed_f == 8'h99; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_153; // @[Reg.scala 27:20]
  wire [1:0] _T_22517 = _T_22056 ? bht_bank_rd_data_out_1_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22772 = _T_22771 | _T_22517; // @[Mux.scala 27:72]
  wire  _T_22059 = bht_rd_addr_hashed_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_154; // @[Reg.scala 27:20]
  wire [1:0] _T_22518 = _T_22059 ? bht_bank_rd_data_out_1_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22773 = _T_22772 | _T_22518; // @[Mux.scala 27:72]
  wire  _T_22062 = bht_rd_addr_hashed_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_155; // @[Reg.scala 27:20]
  wire [1:0] _T_22519 = _T_22062 ? bht_bank_rd_data_out_1_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22774 = _T_22773 | _T_22519; // @[Mux.scala 27:72]
  wire  _T_22065 = bht_rd_addr_hashed_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_156; // @[Reg.scala 27:20]
  wire [1:0] _T_22520 = _T_22065 ? bht_bank_rd_data_out_1_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22775 = _T_22774 | _T_22520; // @[Mux.scala 27:72]
  wire  _T_22068 = bht_rd_addr_hashed_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_157; // @[Reg.scala 27:20]
  wire [1:0] _T_22521 = _T_22068 ? bht_bank_rd_data_out_1_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22776 = _T_22775 | _T_22521; // @[Mux.scala 27:72]
  wire  _T_22071 = bht_rd_addr_hashed_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_158; // @[Reg.scala 27:20]
  wire [1:0] _T_22522 = _T_22071 ? bht_bank_rd_data_out_1_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22777 = _T_22776 | _T_22522; // @[Mux.scala 27:72]
  wire  _T_22074 = bht_rd_addr_hashed_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_159; // @[Reg.scala 27:20]
  wire [1:0] _T_22523 = _T_22074 ? bht_bank_rd_data_out_1_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22778 = _T_22777 | _T_22523; // @[Mux.scala 27:72]
  wire  _T_22077 = bht_rd_addr_hashed_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_160; // @[Reg.scala 27:20]
  wire [1:0] _T_22524 = _T_22077 ? bht_bank_rd_data_out_1_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22779 = _T_22778 | _T_22524; // @[Mux.scala 27:72]
  wire  _T_22080 = bht_rd_addr_hashed_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_161; // @[Reg.scala 27:20]
  wire [1:0] _T_22525 = _T_22080 ? bht_bank_rd_data_out_1_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22780 = _T_22779 | _T_22525; // @[Mux.scala 27:72]
  wire  _T_22083 = bht_rd_addr_hashed_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_162; // @[Reg.scala 27:20]
  wire [1:0] _T_22526 = _T_22083 ? bht_bank_rd_data_out_1_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22781 = _T_22780 | _T_22526; // @[Mux.scala 27:72]
  wire  _T_22086 = bht_rd_addr_hashed_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_163; // @[Reg.scala 27:20]
  wire [1:0] _T_22527 = _T_22086 ? bht_bank_rd_data_out_1_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22782 = _T_22781 | _T_22527; // @[Mux.scala 27:72]
  wire  _T_22089 = bht_rd_addr_hashed_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_164; // @[Reg.scala 27:20]
  wire [1:0] _T_22528 = _T_22089 ? bht_bank_rd_data_out_1_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22783 = _T_22782 | _T_22528; // @[Mux.scala 27:72]
  wire  _T_22092 = bht_rd_addr_hashed_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_165; // @[Reg.scala 27:20]
  wire [1:0] _T_22529 = _T_22092 ? bht_bank_rd_data_out_1_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22784 = _T_22783 | _T_22529; // @[Mux.scala 27:72]
  wire  _T_22095 = bht_rd_addr_hashed_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_166; // @[Reg.scala 27:20]
  wire [1:0] _T_22530 = _T_22095 ? bht_bank_rd_data_out_1_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22785 = _T_22784 | _T_22530; // @[Mux.scala 27:72]
  wire  _T_22098 = bht_rd_addr_hashed_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_167; // @[Reg.scala 27:20]
  wire [1:0] _T_22531 = _T_22098 ? bht_bank_rd_data_out_1_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22786 = _T_22785 | _T_22531; // @[Mux.scala 27:72]
  wire  _T_22101 = bht_rd_addr_hashed_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_168; // @[Reg.scala 27:20]
  wire [1:0] _T_22532 = _T_22101 ? bht_bank_rd_data_out_1_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22787 = _T_22786 | _T_22532; // @[Mux.scala 27:72]
  wire  _T_22104 = bht_rd_addr_hashed_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_169; // @[Reg.scala 27:20]
  wire [1:0] _T_22533 = _T_22104 ? bht_bank_rd_data_out_1_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22788 = _T_22787 | _T_22533; // @[Mux.scala 27:72]
  wire  _T_22107 = bht_rd_addr_hashed_f == 8'haa; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_170; // @[Reg.scala 27:20]
  wire [1:0] _T_22534 = _T_22107 ? bht_bank_rd_data_out_1_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22789 = _T_22788 | _T_22534; // @[Mux.scala 27:72]
  wire  _T_22110 = bht_rd_addr_hashed_f == 8'hab; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_171; // @[Reg.scala 27:20]
  wire [1:0] _T_22535 = _T_22110 ? bht_bank_rd_data_out_1_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22790 = _T_22789 | _T_22535; // @[Mux.scala 27:72]
  wire  _T_22113 = bht_rd_addr_hashed_f == 8'hac; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_172; // @[Reg.scala 27:20]
  wire [1:0] _T_22536 = _T_22113 ? bht_bank_rd_data_out_1_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22791 = _T_22790 | _T_22536; // @[Mux.scala 27:72]
  wire  _T_22116 = bht_rd_addr_hashed_f == 8'had; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_173; // @[Reg.scala 27:20]
  wire [1:0] _T_22537 = _T_22116 ? bht_bank_rd_data_out_1_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22792 = _T_22791 | _T_22537; // @[Mux.scala 27:72]
  wire  _T_22119 = bht_rd_addr_hashed_f == 8'hae; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_174; // @[Reg.scala 27:20]
  wire [1:0] _T_22538 = _T_22119 ? bht_bank_rd_data_out_1_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22793 = _T_22792 | _T_22538; // @[Mux.scala 27:72]
  wire  _T_22122 = bht_rd_addr_hashed_f == 8'haf; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_175; // @[Reg.scala 27:20]
  wire [1:0] _T_22539 = _T_22122 ? bht_bank_rd_data_out_1_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22794 = _T_22793 | _T_22539; // @[Mux.scala 27:72]
  wire  _T_22125 = bht_rd_addr_hashed_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_176; // @[Reg.scala 27:20]
  wire [1:0] _T_22540 = _T_22125 ? bht_bank_rd_data_out_1_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22795 = _T_22794 | _T_22540; // @[Mux.scala 27:72]
  wire  _T_22128 = bht_rd_addr_hashed_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_177; // @[Reg.scala 27:20]
  wire [1:0] _T_22541 = _T_22128 ? bht_bank_rd_data_out_1_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22796 = _T_22795 | _T_22541; // @[Mux.scala 27:72]
  wire  _T_22131 = bht_rd_addr_hashed_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_178; // @[Reg.scala 27:20]
  wire [1:0] _T_22542 = _T_22131 ? bht_bank_rd_data_out_1_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22797 = _T_22796 | _T_22542; // @[Mux.scala 27:72]
  wire  _T_22134 = bht_rd_addr_hashed_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_179; // @[Reg.scala 27:20]
  wire [1:0] _T_22543 = _T_22134 ? bht_bank_rd_data_out_1_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22798 = _T_22797 | _T_22543; // @[Mux.scala 27:72]
  wire  _T_22137 = bht_rd_addr_hashed_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_180; // @[Reg.scala 27:20]
  wire [1:0] _T_22544 = _T_22137 ? bht_bank_rd_data_out_1_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22799 = _T_22798 | _T_22544; // @[Mux.scala 27:72]
  wire  _T_22140 = bht_rd_addr_hashed_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_181; // @[Reg.scala 27:20]
  wire [1:0] _T_22545 = _T_22140 ? bht_bank_rd_data_out_1_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22800 = _T_22799 | _T_22545; // @[Mux.scala 27:72]
  wire  _T_22143 = bht_rd_addr_hashed_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_182; // @[Reg.scala 27:20]
  wire [1:0] _T_22546 = _T_22143 ? bht_bank_rd_data_out_1_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22801 = _T_22800 | _T_22546; // @[Mux.scala 27:72]
  wire  _T_22146 = bht_rd_addr_hashed_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_183; // @[Reg.scala 27:20]
  wire [1:0] _T_22547 = _T_22146 ? bht_bank_rd_data_out_1_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22802 = _T_22801 | _T_22547; // @[Mux.scala 27:72]
  wire  _T_22149 = bht_rd_addr_hashed_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_184; // @[Reg.scala 27:20]
  wire [1:0] _T_22548 = _T_22149 ? bht_bank_rd_data_out_1_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22803 = _T_22802 | _T_22548; // @[Mux.scala 27:72]
  wire  _T_22152 = bht_rd_addr_hashed_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_185; // @[Reg.scala 27:20]
  wire [1:0] _T_22549 = _T_22152 ? bht_bank_rd_data_out_1_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22804 = _T_22803 | _T_22549; // @[Mux.scala 27:72]
  wire  _T_22155 = bht_rd_addr_hashed_f == 8'hba; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_186; // @[Reg.scala 27:20]
  wire [1:0] _T_22550 = _T_22155 ? bht_bank_rd_data_out_1_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22805 = _T_22804 | _T_22550; // @[Mux.scala 27:72]
  wire  _T_22158 = bht_rd_addr_hashed_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_187; // @[Reg.scala 27:20]
  wire [1:0] _T_22551 = _T_22158 ? bht_bank_rd_data_out_1_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22806 = _T_22805 | _T_22551; // @[Mux.scala 27:72]
  wire  _T_22161 = bht_rd_addr_hashed_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_188; // @[Reg.scala 27:20]
  wire [1:0] _T_22552 = _T_22161 ? bht_bank_rd_data_out_1_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22807 = _T_22806 | _T_22552; // @[Mux.scala 27:72]
  wire  _T_22164 = bht_rd_addr_hashed_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_189; // @[Reg.scala 27:20]
  wire [1:0] _T_22553 = _T_22164 ? bht_bank_rd_data_out_1_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22808 = _T_22807 | _T_22553; // @[Mux.scala 27:72]
  wire  _T_22167 = bht_rd_addr_hashed_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_190; // @[Reg.scala 27:20]
  wire [1:0] _T_22554 = _T_22167 ? bht_bank_rd_data_out_1_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22809 = _T_22808 | _T_22554; // @[Mux.scala 27:72]
  wire  _T_22170 = bht_rd_addr_hashed_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_191; // @[Reg.scala 27:20]
  wire [1:0] _T_22555 = _T_22170 ? bht_bank_rd_data_out_1_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22810 = _T_22809 | _T_22555; // @[Mux.scala 27:72]
  wire  _T_22173 = bht_rd_addr_hashed_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_192; // @[Reg.scala 27:20]
  wire [1:0] _T_22556 = _T_22173 ? bht_bank_rd_data_out_1_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22811 = _T_22810 | _T_22556; // @[Mux.scala 27:72]
  wire  _T_22176 = bht_rd_addr_hashed_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_193; // @[Reg.scala 27:20]
  wire [1:0] _T_22557 = _T_22176 ? bht_bank_rd_data_out_1_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22812 = _T_22811 | _T_22557; // @[Mux.scala 27:72]
  wire  _T_22179 = bht_rd_addr_hashed_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_194; // @[Reg.scala 27:20]
  wire [1:0] _T_22558 = _T_22179 ? bht_bank_rd_data_out_1_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22813 = _T_22812 | _T_22558; // @[Mux.scala 27:72]
  wire  _T_22182 = bht_rd_addr_hashed_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_195; // @[Reg.scala 27:20]
  wire [1:0] _T_22559 = _T_22182 ? bht_bank_rd_data_out_1_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22814 = _T_22813 | _T_22559; // @[Mux.scala 27:72]
  wire  _T_22185 = bht_rd_addr_hashed_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_196; // @[Reg.scala 27:20]
  wire [1:0] _T_22560 = _T_22185 ? bht_bank_rd_data_out_1_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22815 = _T_22814 | _T_22560; // @[Mux.scala 27:72]
  wire  _T_22188 = bht_rd_addr_hashed_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_197; // @[Reg.scala 27:20]
  wire [1:0] _T_22561 = _T_22188 ? bht_bank_rd_data_out_1_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22816 = _T_22815 | _T_22561; // @[Mux.scala 27:72]
  wire  _T_22191 = bht_rd_addr_hashed_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_198; // @[Reg.scala 27:20]
  wire [1:0] _T_22562 = _T_22191 ? bht_bank_rd_data_out_1_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22817 = _T_22816 | _T_22562; // @[Mux.scala 27:72]
  wire  _T_22194 = bht_rd_addr_hashed_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_199; // @[Reg.scala 27:20]
  wire [1:0] _T_22563 = _T_22194 ? bht_bank_rd_data_out_1_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22818 = _T_22817 | _T_22563; // @[Mux.scala 27:72]
  wire  _T_22197 = bht_rd_addr_hashed_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_200; // @[Reg.scala 27:20]
  wire [1:0] _T_22564 = _T_22197 ? bht_bank_rd_data_out_1_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22819 = _T_22818 | _T_22564; // @[Mux.scala 27:72]
  wire  _T_22200 = bht_rd_addr_hashed_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_201; // @[Reg.scala 27:20]
  wire [1:0] _T_22565 = _T_22200 ? bht_bank_rd_data_out_1_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22820 = _T_22819 | _T_22565; // @[Mux.scala 27:72]
  wire  _T_22203 = bht_rd_addr_hashed_f == 8'hca; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_202; // @[Reg.scala 27:20]
  wire [1:0] _T_22566 = _T_22203 ? bht_bank_rd_data_out_1_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22821 = _T_22820 | _T_22566; // @[Mux.scala 27:72]
  wire  _T_22206 = bht_rd_addr_hashed_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_203; // @[Reg.scala 27:20]
  wire [1:0] _T_22567 = _T_22206 ? bht_bank_rd_data_out_1_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22822 = _T_22821 | _T_22567; // @[Mux.scala 27:72]
  wire  _T_22209 = bht_rd_addr_hashed_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_204; // @[Reg.scala 27:20]
  wire [1:0] _T_22568 = _T_22209 ? bht_bank_rd_data_out_1_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22823 = _T_22822 | _T_22568; // @[Mux.scala 27:72]
  wire  _T_22212 = bht_rd_addr_hashed_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_205; // @[Reg.scala 27:20]
  wire [1:0] _T_22569 = _T_22212 ? bht_bank_rd_data_out_1_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22824 = _T_22823 | _T_22569; // @[Mux.scala 27:72]
  wire  _T_22215 = bht_rd_addr_hashed_f == 8'hce; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_206; // @[Reg.scala 27:20]
  wire [1:0] _T_22570 = _T_22215 ? bht_bank_rd_data_out_1_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22825 = _T_22824 | _T_22570; // @[Mux.scala 27:72]
  wire  _T_22218 = bht_rd_addr_hashed_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_207; // @[Reg.scala 27:20]
  wire [1:0] _T_22571 = _T_22218 ? bht_bank_rd_data_out_1_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22826 = _T_22825 | _T_22571; // @[Mux.scala 27:72]
  wire  _T_22221 = bht_rd_addr_hashed_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_208; // @[Reg.scala 27:20]
  wire [1:0] _T_22572 = _T_22221 ? bht_bank_rd_data_out_1_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22827 = _T_22826 | _T_22572; // @[Mux.scala 27:72]
  wire  _T_22224 = bht_rd_addr_hashed_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_209; // @[Reg.scala 27:20]
  wire [1:0] _T_22573 = _T_22224 ? bht_bank_rd_data_out_1_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22828 = _T_22827 | _T_22573; // @[Mux.scala 27:72]
  wire  _T_22227 = bht_rd_addr_hashed_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_210; // @[Reg.scala 27:20]
  wire [1:0] _T_22574 = _T_22227 ? bht_bank_rd_data_out_1_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22829 = _T_22828 | _T_22574; // @[Mux.scala 27:72]
  wire  _T_22230 = bht_rd_addr_hashed_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_211; // @[Reg.scala 27:20]
  wire [1:0] _T_22575 = _T_22230 ? bht_bank_rd_data_out_1_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22830 = _T_22829 | _T_22575; // @[Mux.scala 27:72]
  wire  _T_22233 = bht_rd_addr_hashed_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_212; // @[Reg.scala 27:20]
  wire [1:0] _T_22576 = _T_22233 ? bht_bank_rd_data_out_1_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22831 = _T_22830 | _T_22576; // @[Mux.scala 27:72]
  wire  _T_22236 = bht_rd_addr_hashed_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_213; // @[Reg.scala 27:20]
  wire [1:0] _T_22577 = _T_22236 ? bht_bank_rd_data_out_1_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22832 = _T_22831 | _T_22577; // @[Mux.scala 27:72]
  wire  _T_22239 = bht_rd_addr_hashed_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_214; // @[Reg.scala 27:20]
  wire [1:0] _T_22578 = _T_22239 ? bht_bank_rd_data_out_1_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22833 = _T_22832 | _T_22578; // @[Mux.scala 27:72]
  wire  _T_22242 = bht_rd_addr_hashed_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_215; // @[Reg.scala 27:20]
  wire [1:0] _T_22579 = _T_22242 ? bht_bank_rd_data_out_1_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22834 = _T_22833 | _T_22579; // @[Mux.scala 27:72]
  wire  _T_22245 = bht_rd_addr_hashed_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_216; // @[Reg.scala 27:20]
  wire [1:0] _T_22580 = _T_22245 ? bht_bank_rd_data_out_1_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22835 = _T_22834 | _T_22580; // @[Mux.scala 27:72]
  wire  _T_22248 = bht_rd_addr_hashed_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_217; // @[Reg.scala 27:20]
  wire [1:0] _T_22581 = _T_22248 ? bht_bank_rd_data_out_1_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22836 = _T_22835 | _T_22581; // @[Mux.scala 27:72]
  wire  _T_22251 = bht_rd_addr_hashed_f == 8'hda; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_218; // @[Reg.scala 27:20]
  wire [1:0] _T_22582 = _T_22251 ? bht_bank_rd_data_out_1_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22837 = _T_22836 | _T_22582; // @[Mux.scala 27:72]
  wire  _T_22254 = bht_rd_addr_hashed_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_219; // @[Reg.scala 27:20]
  wire [1:0] _T_22583 = _T_22254 ? bht_bank_rd_data_out_1_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22838 = _T_22837 | _T_22583; // @[Mux.scala 27:72]
  wire  _T_22257 = bht_rd_addr_hashed_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_220; // @[Reg.scala 27:20]
  wire [1:0] _T_22584 = _T_22257 ? bht_bank_rd_data_out_1_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22839 = _T_22838 | _T_22584; // @[Mux.scala 27:72]
  wire  _T_22260 = bht_rd_addr_hashed_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_221; // @[Reg.scala 27:20]
  wire [1:0] _T_22585 = _T_22260 ? bht_bank_rd_data_out_1_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22840 = _T_22839 | _T_22585; // @[Mux.scala 27:72]
  wire  _T_22263 = bht_rd_addr_hashed_f == 8'hde; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_222; // @[Reg.scala 27:20]
  wire [1:0] _T_22586 = _T_22263 ? bht_bank_rd_data_out_1_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22841 = _T_22840 | _T_22586; // @[Mux.scala 27:72]
  wire  _T_22266 = bht_rd_addr_hashed_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_223; // @[Reg.scala 27:20]
  wire [1:0] _T_22587 = _T_22266 ? bht_bank_rd_data_out_1_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22842 = _T_22841 | _T_22587; // @[Mux.scala 27:72]
  wire  _T_22269 = bht_rd_addr_hashed_f == 8'he0; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_224; // @[Reg.scala 27:20]
  wire [1:0] _T_22588 = _T_22269 ? bht_bank_rd_data_out_1_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22843 = _T_22842 | _T_22588; // @[Mux.scala 27:72]
  wire  _T_22272 = bht_rd_addr_hashed_f == 8'he1; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_225; // @[Reg.scala 27:20]
  wire [1:0] _T_22589 = _T_22272 ? bht_bank_rd_data_out_1_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22844 = _T_22843 | _T_22589; // @[Mux.scala 27:72]
  wire  _T_22275 = bht_rd_addr_hashed_f == 8'he2; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_226; // @[Reg.scala 27:20]
  wire [1:0] _T_22590 = _T_22275 ? bht_bank_rd_data_out_1_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22845 = _T_22844 | _T_22590; // @[Mux.scala 27:72]
  wire  _T_22278 = bht_rd_addr_hashed_f == 8'he3; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_227; // @[Reg.scala 27:20]
  wire [1:0] _T_22591 = _T_22278 ? bht_bank_rd_data_out_1_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22846 = _T_22845 | _T_22591; // @[Mux.scala 27:72]
  wire  _T_22281 = bht_rd_addr_hashed_f == 8'he4; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_228; // @[Reg.scala 27:20]
  wire [1:0] _T_22592 = _T_22281 ? bht_bank_rd_data_out_1_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22847 = _T_22846 | _T_22592; // @[Mux.scala 27:72]
  wire  _T_22284 = bht_rd_addr_hashed_f == 8'he5; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_229; // @[Reg.scala 27:20]
  wire [1:0] _T_22593 = _T_22284 ? bht_bank_rd_data_out_1_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22848 = _T_22847 | _T_22593; // @[Mux.scala 27:72]
  wire  _T_22287 = bht_rd_addr_hashed_f == 8'he6; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_230; // @[Reg.scala 27:20]
  wire [1:0] _T_22594 = _T_22287 ? bht_bank_rd_data_out_1_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22849 = _T_22848 | _T_22594; // @[Mux.scala 27:72]
  wire  _T_22290 = bht_rd_addr_hashed_f == 8'he7; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_231; // @[Reg.scala 27:20]
  wire [1:0] _T_22595 = _T_22290 ? bht_bank_rd_data_out_1_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22850 = _T_22849 | _T_22595; // @[Mux.scala 27:72]
  wire  _T_22293 = bht_rd_addr_hashed_f == 8'he8; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_232; // @[Reg.scala 27:20]
  wire [1:0] _T_22596 = _T_22293 ? bht_bank_rd_data_out_1_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22851 = _T_22850 | _T_22596; // @[Mux.scala 27:72]
  wire  _T_22296 = bht_rd_addr_hashed_f == 8'he9; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_233; // @[Reg.scala 27:20]
  wire [1:0] _T_22597 = _T_22296 ? bht_bank_rd_data_out_1_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22852 = _T_22851 | _T_22597; // @[Mux.scala 27:72]
  wire  _T_22299 = bht_rd_addr_hashed_f == 8'hea; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_234; // @[Reg.scala 27:20]
  wire [1:0] _T_22598 = _T_22299 ? bht_bank_rd_data_out_1_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22853 = _T_22852 | _T_22598; // @[Mux.scala 27:72]
  wire  _T_22302 = bht_rd_addr_hashed_f == 8'heb; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_235; // @[Reg.scala 27:20]
  wire [1:0] _T_22599 = _T_22302 ? bht_bank_rd_data_out_1_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22854 = _T_22853 | _T_22599; // @[Mux.scala 27:72]
  wire  _T_22305 = bht_rd_addr_hashed_f == 8'hec; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_236; // @[Reg.scala 27:20]
  wire [1:0] _T_22600 = _T_22305 ? bht_bank_rd_data_out_1_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22855 = _T_22854 | _T_22600; // @[Mux.scala 27:72]
  wire  _T_22308 = bht_rd_addr_hashed_f == 8'hed; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_237; // @[Reg.scala 27:20]
  wire [1:0] _T_22601 = _T_22308 ? bht_bank_rd_data_out_1_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22856 = _T_22855 | _T_22601; // @[Mux.scala 27:72]
  wire  _T_22311 = bht_rd_addr_hashed_f == 8'hee; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_238; // @[Reg.scala 27:20]
  wire [1:0] _T_22602 = _T_22311 ? bht_bank_rd_data_out_1_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22857 = _T_22856 | _T_22602; // @[Mux.scala 27:72]
  wire  _T_22314 = bht_rd_addr_hashed_f == 8'hef; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_239; // @[Reg.scala 27:20]
  wire [1:0] _T_22603 = _T_22314 ? bht_bank_rd_data_out_1_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22858 = _T_22857 | _T_22603; // @[Mux.scala 27:72]
  wire  _T_22317 = bht_rd_addr_hashed_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_240; // @[Reg.scala 27:20]
  wire [1:0] _T_22604 = _T_22317 ? bht_bank_rd_data_out_1_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22859 = _T_22858 | _T_22604; // @[Mux.scala 27:72]
  wire  _T_22320 = bht_rd_addr_hashed_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_241; // @[Reg.scala 27:20]
  wire [1:0] _T_22605 = _T_22320 ? bht_bank_rd_data_out_1_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22860 = _T_22859 | _T_22605; // @[Mux.scala 27:72]
  wire  _T_22323 = bht_rd_addr_hashed_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_242; // @[Reg.scala 27:20]
  wire [1:0] _T_22606 = _T_22323 ? bht_bank_rd_data_out_1_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22861 = _T_22860 | _T_22606; // @[Mux.scala 27:72]
  wire  _T_22326 = bht_rd_addr_hashed_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_243; // @[Reg.scala 27:20]
  wire [1:0] _T_22607 = _T_22326 ? bht_bank_rd_data_out_1_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22862 = _T_22861 | _T_22607; // @[Mux.scala 27:72]
  wire  _T_22329 = bht_rd_addr_hashed_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_244; // @[Reg.scala 27:20]
  wire [1:0] _T_22608 = _T_22329 ? bht_bank_rd_data_out_1_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22863 = _T_22862 | _T_22608; // @[Mux.scala 27:72]
  wire  _T_22332 = bht_rd_addr_hashed_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_245; // @[Reg.scala 27:20]
  wire [1:0] _T_22609 = _T_22332 ? bht_bank_rd_data_out_1_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22864 = _T_22863 | _T_22609; // @[Mux.scala 27:72]
  wire  _T_22335 = bht_rd_addr_hashed_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_246; // @[Reg.scala 27:20]
  wire [1:0] _T_22610 = _T_22335 ? bht_bank_rd_data_out_1_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22865 = _T_22864 | _T_22610; // @[Mux.scala 27:72]
  wire  _T_22338 = bht_rd_addr_hashed_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_247; // @[Reg.scala 27:20]
  wire [1:0] _T_22611 = _T_22338 ? bht_bank_rd_data_out_1_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22866 = _T_22865 | _T_22611; // @[Mux.scala 27:72]
  wire  _T_22341 = bht_rd_addr_hashed_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_248; // @[Reg.scala 27:20]
  wire [1:0] _T_22612 = _T_22341 ? bht_bank_rd_data_out_1_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22867 = _T_22866 | _T_22612; // @[Mux.scala 27:72]
  wire  _T_22344 = bht_rd_addr_hashed_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_249; // @[Reg.scala 27:20]
  wire [1:0] _T_22613 = _T_22344 ? bht_bank_rd_data_out_1_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22868 = _T_22867 | _T_22613; // @[Mux.scala 27:72]
  wire  _T_22347 = bht_rd_addr_hashed_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_250; // @[Reg.scala 27:20]
  wire [1:0] _T_22614 = _T_22347 ? bht_bank_rd_data_out_1_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22869 = _T_22868 | _T_22614; // @[Mux.scala 27:72]
  wire  _T_22350 = bht_rd_addr_hashed_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_251; // @[Reg.scala 27:20]
  wire [1:0] _T_22615 = _T_22350 ? bht_bank_rd_data_out_1_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22870 = _T_22869 | _T_22615; // @[Mux.scala 27:72]
  wire  _T_22353 = bht_rd_addr_hashed_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_252; // @[Reg.scala 27:20]
  wire [1:0] _T_22616 = _T_22353 ? bht_bank_rd_data_out_1_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22871 = _T_22870 | _T_22616; // @[Mux.scala 27:72]
  wire  _T_22356 = bht_rd_addr_hashed_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_253; // @[Reg.scala 27:20]
  wire [1:0] _T_22617 = _T_22356 ? bht_bank_rd_data_out_1_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22872 = _T_22871 | _T_22617; // @[Mux.scala 27:72]
  wire  _T_22359 = bht_rd_addr_hashed_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_254; // @[Reg.scala 27:20]
  wire [1:0] _T_22618 = _T_22359 ? bht_bank_rd_data_out_1_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22873 = _T_22872 | _T_22618; // @[Mux.scala 27:72]
  wire  _T_22362 = bht_rd_addr_hashed_f == 8'hff; // @[el2_ifu_bp_ctl.scala 396:106]
  reg [1:0] bht_bank_rd_data_out_1_255; // @[Reg.scala 27:20]
  wire [1:0] _T_22619 = _T_22362 ? bht_bank_rd_data_out_1_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank1_rd_data_f = _T_22873 | _T_22619; // @[Mux.scala 27:72]
  wire [1:0] _T_258 = _T_143 ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [9:0] _T_569 = {btb_rd_addr_p1_f,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_rd_addr_hashed_p1_f = _T_569[9:2] ^ fghr; // @[el2_lib.scala 191:35]
  wire  _T_22877 = bht_rd_addr_hashed_p1_f == 8'h0; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23644 = _T_22877 ? bht_bank_rd_data_out_1_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_22880 = bht_rd_addr_hashed_p1_f == 8'h1; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23645 = _T_22880 ? bht_bank_rd_data_out_1_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23900 = _T_23644 | _T_23645; // @[Mux.scala 27:72]
  wire  _T_22883 = bht_rd_addr_hashed_p1_f == 8'h2; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23646 = _T_22883 ? bht_bank_rd_data_out_1_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23901 = _T_23900 | _T_23646; // @[Mux.scala 27:72]
  wire  _T_22886 = bht_rd_addr_hashed_p1_f == 8'h3; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23647 = _T_22886 ? bht_bank_rd_data_out_1_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23902 = _T_23901 | _T_23647; // @[Mux.scala 27:72]
  wire  _T_22889 = bht_rd_addr_hashed_p1_f == 8'h4; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23648 = _T_22889 ? bht_bank_rd_data_out_1_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23903 = _T_23902 | _T_23648; // @[Mux.scala 27:72]
  wire  _T_22892 = bht_rd_addr_hashed_p1_f == 8'h5; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23649 = _T_22892 ? bht_bank_rd_data_out_1_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23904 = _T_23903 | _T_23649; // @[Mux.scala 27:72]
  wire  _T_22895 = bht_rd_addr_hashed_p1_f == 8'h6; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23650 = _T_22895 ? bht_bank_rd_data_out_1_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23905 = _T_23904 | _T_23650; // @[Mux.scala 27:72]
  wire  _T_22898 = bht_rd_addr_hashed_p1_f == 8'h7; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23651 = _T_22898 ? bht_bank_rd_data_out_1_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23906 = _T_23905 | _T_23651; // @[Mux.scala 27:72]
  wire  _T_22901 = bht_rd_addr_hashed_p1_f == 8'h8; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23652 = _T_22901 ? bht_bank_rd_data_out_1_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23907 = _T_23906 | _T_23652; // @[Mux.scala 27:72]
  wire  _T_22904 = bht_rd_addr_hashed_p1_f == 8'h9; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23653 = _T_22904 ? bht_bank_rd_data_out_1_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23908 = _T_23907 | _T_23653; // @[Mux.scala 27:72]
  wire  _T_22907 = bht_rd_addr_hashed_p1_f == 8'ha; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23654 = _T_22907 ? bht_bank_rd_data_out_1_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23909 = _T_23908 | _T_23654; // @[Mux.scala 27:72]
  wire  _T_22910 = bht_rd_addr_hashed_p1_f == 8'hb; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23655 = _T_22910 ? bht_bank_rd_data_out_1_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23910 = _T_23909 | _T_23655; // @[Mux.scala 27:72]
  wire  _T_22913 = bht_rd_addr_hashed_p1_f == 8'hc; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23656 = _T_22913 ? bht_bank_rd_data_out_1_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23911 = _T_23910 | _T_23656; // @[Mux.scala 27:72]
  wire  _T_22916 = bht_rd_addr_hashed_p1_f == 8'hd; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23657 = _T_22916 ? bht_bank_rd_data_out_1_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23912 = _T_23911 | _T_23657; // @[Mux.scala 27:72]
  wire  _T_22919 = bht_rd_addr_hashed_p1_f == 8'he; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23658 = _T_22919 ? bht_bank_rd_data_out_1_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23913 = _T_23912 | _T_23658; // @[Mux.scala 27:72]
  wire  _T_22922 = bht_rd_addr_hashed_p1_f == 8'hf; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23659 = _T_22922 ? bht_bank_rd_data_out_1_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23914 = _T_23913 | _T_23659; // @[Mux.scala 27:72]
  wire  _T_22925 = bht_rd_addr_hashed_p1_f == 8'h10; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23660 = _T_22925 ? bht_bank_rd_data_out_1_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23915 = _T_23914 | _T_23660; // @[Mux.scala 27:72]
  wire  _T_22928 = bht_rd_addr_hashed_p1_f == 8'h11; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23661 = _T_22928 ? bht_bank_rd_data_out_1_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23916 = _T_23915 | _T_23661; // @[Mux.scala 27:72]
  wire  _T_22931 = bht_rd_addr_hashed_p1_f == 8'h12; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23662 = _T_22931 ? bht_bank_rd_data_out_1_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23917 = _T_23916 | _T_23662; // @[Mux.scala 27:72]
  wire  _T_22934 = bht_rd_addr_hashed_p1_f == 8'h13; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23663 = _T_22934 ? bht_bank_rd_data_out_1_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23918 = _T_23917 | _T_23663; // @[Mux.scala 27:72]
  wire  _T_22937 = bht_rd_addr_hashed_p1_f == 8'h14; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23664 = _T_22937 ? bht_bank_rd_data_out_1_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23919 = _T_23918 | _T_23664; // @[Mux.scala 27:72]
  wire  _T_22940 = bht_rd_addr_hashed_p1_f == 8'h15; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23665 = _T_22940 ? bht_bank_rd_data_out_1_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23920 = _T_23919 | _T_23665; // @[Mux.scala 27:72]
  wire  _T_22943 = bht_rd_addr_hashed_p1_f == 8'h16; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23666 = _T_22943 ? bht_bank_rd_data_out_1_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23921 = _T_23920 | _T_23666; // @[Mux.scala 27:72]
  wire  _T_22946 = bht_rd_addr_hashed_p1_f == 8'h17; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23667 = _T_22946 ? bht_bank_rd_data_out_1_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23922 = _T_23921 | _T_23667; // @[Mux.scala 27:72]
  wire  _T_22949 = bht_rd_addr_hashed_p1_f == 8'h18; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23668 = _T_22949 ? bht_bank_rd_data_out_1_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23923 = _T_23922 | _T_23668; // @[Mux.scala 27:72]
  wire  _T_22952 = bht_rd_addr_hashed_p1_f == 8'h19; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23669 = _T_22952 ? bht_bank_rd_data_out_1_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23924 = _T_23923 | _T_23669; // @[Mux.scala 27:72]
  wire  _T_22955 = bht_rd_addr_hashed_p1_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23670 = _T_22955 ? bht_bank_rd_data_out_1_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23925 = _T_23924 | _T_23670; // @[Mux.scala 27:72]
  wire  _T_22958 = bht_rd_addr_hashed_p1_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23671 = _T_22958 ? bht_bank_rd_data_out_1_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23926 = _T_23925 | _T_23671; // @[Mux.scala 27:72]
  wire  _T_22961 = bht_rd_addr_hashed_p1_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23672 = _T_22961 ? bht_bank_rd_data_out_1_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23927 = _T_23926 | _T_23672; // @[Mux.scala 27:72]
  wire  _T_22964 = bht_rd_addr_hashed_p1_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23673 = _T_22964 ? bht_bank_rd_data_out_1_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23928 = _T_23927 | _T_23673; // @[Mux.scala 27:72]
  wire  _T_22967 = bht_rd_addr_hashed_p1_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23674 = _T_22967 ? bht_bank_rd_data_out_1_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23929 = _T_23928 | _T_23674; // @[Mux.scala 27:72]
  wire  _T_22970 = bht_rd_addr_hashed_p1_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23675 = _T_22970 ? bht_bank_rd_data_out_1_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23930 = _T_23929 | _T_23675; // @[Mux.scala 27:72]
  wire  _T_22973 = bht_rd_addr_hashed_p1_f == 8'h20; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23676 = _T_22973 ? bht_bank_rd_data_out_1_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23931 = _T_23930 | _T_23676; // @[Mux.scala 27:72]
  wire  _T_22976 = bht_rd_addr_hashed_p1_f == 8'h21; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23677 = _T_22976 ? bht_bank_rd_data_out_1_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23932 = _T_23931 | _T_23677; // @[Mux.scala 27:72]
  wire  _T_22979 = bht_rd_addr_hashed_p1_f == 8'h22; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23678 = _T_22979 ? bht_bank_rd_data_out_1_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23933 = _T_23932 | _T_23678; // @[Mux.scala 27:72]
  wire  _T_22982 = bht_rd_addr_hashed_p1_f == 8'h23; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23679 = _T_22982 ? bht_bank_rd_data_out_1_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23934 = _T_23933 | _T_23679; // @[Mux.scala 27:72]
  wire  _T_22985 = bht_rd_addr_hashed_p1_f == 8'h24; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23680 = _T_22985 ? bht_bank_rd_data_out_1_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23935 = _T_23934 | _T_23680; // @[Mux.scala 27:72]
  wire  _T_22988 = bht_rd_addr_hashed_p1_f == 8'h25; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23681 = _T_22988 ? bht_bank_rd_data_out_1_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23936 = _T_23935 | _T_23681; // @[Mux.scala 27:72]
  wire  _T_22991 = bht_rd_addr_hashed_p1_f == 8'h26; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23682 = _T_22991 ? bht_bank_rd_data_out_1_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23937 = _T_23936 | _T_23682; // @[Mux.scala 27:72]
  wire  _T_22994 = bht_rd_addr_hashed_p1_f == 8'h27; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23683 = _T_22994 ? bht_bank_rd_data_out_1_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23938 = _T_23937 | _T_23683; // @[Mux.scala 27:72]
  wire  _T_22997 = bht_rd_addr_hashed_p1_f == 8'h28; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23684 = _T_22997 ? bht_bank_rd_data_out_1_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23939 = _T_23938 | _T_23684; // @[Mux.scala 27:72]
  wire  _T_23000 = bht_rd_addr_hashed_p1_f == 8'h29; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23685 = _T_23000 ? bht_bank_rd_data_out_1_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23940 = _T_23939 | _T_23685; // @[Mux.scala 27:72]
  wire  _T_23003 = bht_rd_addr_hashed_p1_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23686 = _T_23003 ? bht_bank_rd_data_out_1_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23941 = _T_23940 | _T_23686; // @[Mux.scala 27:72]
  wire  _T_23006 = bht_rd_addr_hashed_p1_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23687 = _T_23006 ? bht_bank_rd_data_out_1_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23942 = _T_23941 | _T_23687; // @[Mux.scala 27:72]
  wire  _T_23009 = bht_rd_addr_hashed_p1_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23688 = _T_23009 ? bht_bank_rd_data_out_1_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23943 = _T_23942 | _T_23688; // @[Mux.scala 27:72]
  wire  _T_23012 = bht_rd_addr_hashed_p1_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23689 = _T_23012 ? bht_bank_rd_data_out_1_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23944 = _T_23943 | _T_23689; // @[Mux.scala 27:72]
  wire  _T_23015 = bht_rd_addr_hashed_p1_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23690 = _T_23015 ? bht_bank_rd_data_out_1_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23945 = _T_23944 | _T_23690; // @[Mux.scala 27:72]
  wire  _T_23018 = bht_rd_addr_hashed_p1_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23691 = _T_23018 ? bht_bank_rd_data_out_1_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23946 = _T_23945 | _T_23691; // @[Mux.scala 27:72]
  wire  _T_23021 = bht_rd_addr_hashed_p1_f == 8'h30; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23692 = _T_23021 ? bht_bank_rd_data_out_1_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23947 = _T_23946 | _T_23692; // @[Mux.scala 27:72]
  wire  _T_23024 = bht_rd_addr_hashed_p1_f == 8'h31; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23693 = _T_23024 ? bht_bank_rd_data_out_1_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23948 = _T_23947 | _T_23693; // @[Mux.scala 27:72]
  wire  _T_23027 = bht_rd_addr_hashed_p1_f == 8'h32; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23694 = _T_23027 ? bht_bank_rd_data_out_1_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23949 = _T_23948 | _T_23694; // @[Mux.scala 27:72]
  wire  _T_23030 = bht_rd_addr_hashed_p1_f == 8'h33; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23695 = _T_23030 ? bht_bank_rd_data_out_1_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23950 = _T_23949 | _T_23695; // @[Mux.scala 27:72]
  wire  _T_23033 = bht_rd_addr_hashed_p1_f == 8'h34; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23696 = _T_23033 ? bht_bank_rd_data_out_1_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23951 = _T_23950 | _T_23696; // @[Mux.scala 27:72]
  wire  _T_23036 = bht_rd_addr_hashed_p1_f == 8'h35; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23697 = _T_23036 ? bht_bank_rd_data_out_1_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23952 = _T_23951 | _T_23697; // @[Mux.scala 27:72]
  wire  _T_23039 = bht_rd_addr_hashed_p1_f == 8'h36; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23698 = _T_23039 ? bht_bank_rd_data_out_1_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23953 = _T_23952 | _T_23698; // @[Mux.scala 27:72]
  wire  _T_23042 = bht_rd_addr_hashed_p1_f == 8'h37; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23699 = _T_23042 ? bht_bank_rd_data_out_1_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23954 = _T_23953 | _T_23699; // @[Mux.scala 27:72]
  wire  _T_23045 = bht_rd_addr_hashed_p1_f == 8'h38; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23700 = _T_23045 ? bht_bank_rd_data_out_1_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23955 = _T_23954 | _T_23700; // @[Mux.scala 27:72]
  wire  _T_23048 = bht_rd_addr_hashed_p1_f == 8'h39; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23701 = _T_23048 ? bht_bank_rd_data_out_1_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23956 = _T_23955 | _T_23701; // @[Mux.scala 27:72]
  wire  _T_23051 = bht_rd_addr_hashed_p1_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23702 = _T_23051 ? bht_bank_rd_data_out_1_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23957 = _T_23956 | _T_23702; // @[Mux.scala 27:72]
  wire  _T_23054 = bht_rd_addr_hashed_p1_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23703 = _T_23054 ? bht_bank_rd_data_out_1_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23958 = _T_23957 | _T_23703; // @[Mux.scala 27:72]
  wire  _T_23057 = bht_rd_addr_hashed_p1_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23704 = _T_23057 ? bht_bank_rd_data_out_1_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23959 = _T_23958 | _T_23704; // @[Mux.scala 27:72]
  wire  _T_23060 = bht_rd_addr_hashed_p1_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23705 = _T_23060 ? bht_bank_rd_data_out_1_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23960 = _T_23959 | _T_23705; // @[Mux.scala 27:72]
  wire  _T_23063 = bht_rd_addr_hashed_p1_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23706 = _T_23063 ? bht_bank_rd_data_out_1_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23961 = _T_23960 | _T_23706; // @[Mux.scala 27:72]
  wire  _T_23066 = bht_rd_addr_hashed_p1_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23707 = _T_23066 ? bht_bank_rd_data_out_1_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23962 = _T_23961 | _T_23707; // @[Mux.scala 27:72]
  wire  _T_23069 = bht_rd_addr_hashed_p1_f == 8'h40; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23708 = _T_23069 ? bht_bank_rd_data_out_1_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23963 = _T_23962 | _T_23708; // @[Mux.scala 27:72]
  wire  _T_23072 = bht_rd_addr_hashed_p1_f == 8'h41; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23709 = _T_23072 ? bht_bank_rd_data_out_1_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23964 = _T_23963 | _T_23709; // @[Mux.scala 27:72]
  wire  _T_23075 = bht_rd_addr_hashed_p1_f == 8'h42; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23710 = _T_23075 ? bht_bank_rd_data_out_1_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23965 = _T_23964 | _T_23710; // @[Mux.scala 27:72]
  wire  _T_23078 = bht_rd_addr_hashed_p1_f == 8'h43; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23711 = _T_23078 ? bht_bank_rd_data_out_1_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23966 = _T_23965 | _T_23711; // @[Mux.scala 27:72]
  wire  _T_23081 = bht_rd_addr_hashed_p1_f == 8'h44; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23712 = _T_23081 ? bht_bank_rd_data_out_1_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23967 = _T_23966 | _T_23712; // @[Mux.scala 27:72]
  wire  _T_23084 = bht_rd_addr_hashed_p1_f == 8'h45; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23713 = _T_23084 ? bht_bank_rd_data_out_1_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23968 = _T_23967 | _T_23713; // @[Mux.scala 27:72]
  wire  _T_23087 = bht_rd_addr_hashed_p1_f == 8'h46; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23714 = _T_23087 ? bht_bank_rd_data_out_1_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23969 = _T_23968 | _T_23714; // @[Mux.scala 27:72]
  wire  _T_23090 = bht_rd_addr_hashed_p1_f == 8'h47; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23715 = _T_23090 ? bht_bank_rd_data_out_1_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23970 = _T_23969 | _T_23715; // @[Mux.scala 27:72]
  wire  _T_23093 = bht_rd_addr_hashed_p1_f == 8'h48; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23716 = _T_23093 ? bht_bank_rd_data_out_1_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23971 = _T_23970 | _T_23716; // @[Mux.scala 27:72]
  wire  _T_23096 = bht_rd_addr_hashed_p1_f == 8'h49; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23717 = _T_23096 ? bht_bank_rd_data_out_1_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23972 = _T_23971 | _T_23717; // @[Mux.scala 27:72]
  wire  _T_23099 = bht_rd_addr_hashed_p1_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23718 = _T_23099 ? bht_bank_rd_data_out_1_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23973 = _T_23972 | _T_23718; // @[Mux.scala 27:72]
  wire  _T_23102 = bht_rd_addr_hashed_p1_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23719 = _T_23102 ? bht_bank_rd_data_out_1_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23974 = _T_23973 | _T_23719; // @[Mux.scala 27:72]
  wire  _T_23105 = bht_rd_addr_hashed_p1_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23720 = _T_23105 ? bht_bank_rd_data_out_1_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23975 = _T_23974 | _T_23720; // @[Mux.scala 27:72]
  wire  _T_23108 = bht_rd_addr_hashed_p1_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23721 = _T_23108 ? bht_bank_rd_data_out_1_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23976 = _T_23975 | _T_23721; // @[Mux.scala 27:72]
  wire  _T_23111 = bht_rd_addr_hashed_p1_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23722 = _T_23111 ? bht_bank_rd_data_out_1_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23977 = _T_23976 | _T_23722; // @[Mux.scala 27:72]
  wire  _T_23114 = bht_rd_addr_hashed_p1_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23723 = _T_23114 ? bht_bank_rd_data_out_1_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23978 = _T_23977 | _T_23723; // @[Mux.scala 27:72]
  wire  _T_23117 = bht_rd_addr_hashed_p1_f == 8'h50; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23724 = _T_23117 ? bht_bank_rd_data_out_1_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23979 = _T_23978 | _T_23724; // @[Mux.scala 27:72]
  wire  _T_23120 = bht_rd_addr_hashed_p1_f == 8'h51; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23725 = _T_23120 ? bht_bank_rd_data_out_1_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23980 = _T_23979 | _T_23725; // @[Mux.scala 27:72]
  wire  _T_23123 = bht_rd_addr_hashed_p1_f == 8'h52; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23726 = _T_23123 ? bht_bank_rd_data_out_1_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23981 = _T_23980 | _T_23726; // @[Mux.scala 27:72]
  wire  _T_23126 = bht_rd_addr_hashed_p1_f == 8'h53; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23727 = _T_23126 ? bht_bank_rd_data_out_1_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23982 = _T_23981 | _T_23727; // @[Mux.scala 27:72]
  wire  _T_23129 = bht_rd_addr_hashed_p1_f == 8'h54; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23728 = _T_23129 ? bht_bank_rd_data_out_1_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23983 = _T_23982 | _T_23728; // @[Mux.scala 27:72]
  wire  _T_23132 = bht_rd_addr_hashed_p1_f == 8'h55; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23729 = _T_23132 ? bht_bank_rd_data_out_1_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23984 = _T_23983 | _T_23729; // @[Mux.scala 27:72]
  wire  _T_23135 = bht_rd_addr_hashed_p1_f == 8'h56; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23730 = _T_23135 ? bht_bank_rd_data_out_1_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23985 = _T_23984 | _T_23730; // @[Mux.scala 27:72]
  wire  _T_23138 = bht_rd_addr_hashed_p1_f == 8'h57; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23731 = _T_23138 ? bht_bank_rd_data_out_1_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23986 = _T_23985 | _T_23731; // @[Mux.scala 27:72]
  wire  _T_23141 = bht_rd_addr_hashed_p1_f == 8'h58; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23732 = _T_23141 ? bht_bank_rd_data_out_1_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23987 = _T_23986 | _T_23732; // @[Mux.scala 27:72]
  wire  _T_23144 = bht_rd_addr_hashed_p1_f == 8'h59; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23733 = _T_23144 ? bht_bank_rd_data_out_1_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23988 = _T_23987 | _T_23733; // @[Mux.scala 27:72]
  wire  _T_23147 = bht_rd_addr_hashed_p1_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23734 = _T_23147 ? bht_bank_rd_data_out_1_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23989 = _T_23988 | _T_23734; // @[Mux.scala 27:72]
  wire  _T_23150 = bht_rd_addr_hashed_p1_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23735 = _T_23150 ? bht_bank_rd_data_out_1_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23990 = _T_23989 | _T_23735; // @[Mux.scala 27:72]
  wire  _T_23153 = bht_rd_addr_hashed_p1_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23736 = _T_23153 ? bht_bank_rd_data_out_1_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23991 = _T_23990 | _T_23736; // @[Mux.scala 27:72]
  wire  _T_23156 = bht_rd_addr_hashed_p1_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23737 = _T_23156 ? bht_bank_rd_data_out_1_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23992 = _T_23991 | _T_23737; // @[Mux.scala 27:72]
  wire  _T_23159 = bht_rd_addr_hashed_p1_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23738 = _T_23159 ? bht_bank_rd_data_out_1_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23993 = _T_23992 | _T_23738; // @[Mux.scala 27:72]
  wire  _T_23162 = bht_rd_addr_hashed_p1_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23739 = _T_23162 ? bht_bank_rd_data_out_1_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23994 = _T_23993 | _T_23739; // @[Mux.scala 27:72]
  wire  _T_23165 = bht_rd_addr_hashed_p1_f == 8'h60; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23740 = _T_23165 ? bht_bank_rd_data_out_1_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23995 = _T_23994 | _T_23740; // @[Mux.scala 27:72]
  wire  _T_23168 = bht_rd_addr_hashed_p1_f == 8'h61; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23741 = _T_23168 ? bht_bank_rd_data_out_1_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23996 = _T_23995 | _T_23741; // @[Mux.scala 27:72]
  wire  _T_23171 = bht_rd_addr_hashed_p1_f == 8'h62; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23742 = _T_23171 ? bht_bank_rd_data_out_1_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23997 = _T_23996 | _T_23742; // @[Mux.scala 27:72]
  wire  _T_23174 = bht_rd_addr_hashed_p1_f == 8'h63; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23743 = _T_23174 ? bht_bank_rd_data_out_1_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23998 = _T_23997 | _T_23743; // @[Mux.scala 27:72]
  wire  _T_23177 = bht_rd_addr_hashed_p1_f == 8'h64; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23744 = _T_23177 ? bht_bank_rd_data_out_1_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23999 = _T_23998 | _T_23744; // @[Mux.scala 27:72]
  wire  _T_23180 = bht_rd_addr_hashed_p1_f == 8'h65; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23745 = _T_23180 ? bht_bank_rd_data_out_1_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24000 = _T_23999 | _T_23745; // @[Mux.scala 27:72]
  wire  _T_23183 = bht_rd_addr_hashed_p1_f == 8'h66; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23746 = _T_23183 ? bht_bank_rd_data_out_1_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24001 = _T_24000 | _T_23746; // @[Mux.scala 27:72]
  wire  _T_23186 = bht_rd_addr_hashed_p1_f == 8'h67; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23747 = _T_23186 ? bht_bank_rd_data_out_1_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24002 = _T_24001 | _T_23747; // @[Mux.scala 27:72]
  wire  _T_23189 = bht_rd_addr_hashed_p1_f == 8'h68; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23748 = _T_23189 ? bht_bank_rd_data_out_1_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24003 = _T_24002 | _T_23748; // @[Mux.scala 27:72]
  wire  _T_23192 = bht_rd_addr_hashed_p1_f == 8'h69; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23749 = _T_23192 ? bht_bank_rd_data_out_1_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24004 = _T_24003 | _T_23749; // @[Mux.scala 27:72]
  wire  _T_23195 = bht_rd_addr_hashed_p1_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23750 = _T_23195 ? bht_bank_rd_data_out_1_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24005 = _T_24004 | _T_23750; // @[Mux.scala 27:72]
  wire  _T_23198 = bht_rd_addr_hashed_p1_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23751 = _T_23198 ? bht_bank_rd_data_out_1_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24006 = _T_24005 | _T_23751; // @[Mux.scala 27:72]
  wire  _T_23201 = bht_rd_addr_hashed_p1_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23752 = _T_23201 ? bht_bank_rd_data_out_1_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24007 = _T_24006 | _T_23752; // @[Mux.scala 27:72]
  wire  _T_23204 = bht_rd_addr_hashed_p1_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23753 = _T_23204 ? bht_bank_rd_data_out_1_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24008 = _T_24007 | _T_23753; // @[Mux.scala 27:72]
  wire  _T_23207 = bht_rd_addr_hashed_p1_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23754 = _T_23207 ? bht_bank_rd_data_out_1_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24009 = _T_24008 | _T_23754; // @[Mux.scala 27:72]
  wire  _T_23210 = bht_rd_addr_hashed_p1_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23755 = _T_23210 ? bht_bank_rd_data_out_1_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24010 = _T_24009 | _T_23755; // @[Mux.scala 27:72]
  wire  _T_23213 = bht_rd_addr_hashed_p1_f == 8'h70; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23756 = _T_23213 ? bht_bank_rd_data_out_1_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24011 = _T_24010 | _T_23756; // @[Mux.scala 27:72]
  wire  _T_23216 = bht_rd_addr_hashed_p1_f == 8'h71; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23757 = _T_23216 ? bht_bank_rd_data_out_1_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24012 = _T_24011 | _T_23757; // @[Mux.scala 27:72]
  wire  _T_23219 = bht_rd_addr_hashed_p1_f == 8'h72; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23758 = _T_23219 ? bht_bank_rd_data_out_1_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24013 = _T_24012 | _T_23758; // @[Mux.scala 27:72]
  wire  _T_23222 = bht_rd_addr_hashed_p1_f == 8'h73; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23759 = _T_23222 ? bht_bank_rd_data_out_1_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24014 = _T_24013 | _T_23759; // @[Mux.scala 27:72]
  wire  _T_23225 = bht_rd_addr_hashed_p1_f == 8'h74; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23760 = _T_23225 ? bht_bank_rd_data_out_1_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24015 = _T_24014 | _T_23760; // @[Mux.scala 27:72]
  wire  _T_23228 = bht_rd_addr_hashed_p1_f == 8'h75; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23761 = _T_23228 ? bht_bank_rd_data_out_1_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24016 = _T_24015 | _T_23761; // @[Mux.scala 27:72]
  wire  _T_23231 = bht_rd_addr_hashed_p1_f == 8'h76; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23762 = _T_23231 ? bht_bank_rd_data_out_1_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24017 = _T_24016 | _T_23762; // @[Mux.scala 27:72]
  wire  _T_23234 = bht_rd_addr_hashed_p1_f == 8'h77; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23763 = _T_23234 ? bht_bank_rd_data_out_1_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24018 = _T_24017 | _T_23763; // @[Mux.scala 27:72]
  wire  _T_23237 = bht_rd_addr_hashed_p1_f == 8'h78; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23764 = _T_23237 ? bht_bank_rd_data_out_1_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24019 = _T_24018 | _T_23764; // @[Mux.scala 27:72]
  wire  _T_23240 = bht_rd_addr_hashed_p1_f == 8'h79; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23765 = _T_23240 ? bht_bank_rd_data_out_1_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24020 = _T_24019 | _T_23765; // @[Mux.scala 27:72]
  wire  _T_23243 = bht_rd_addr_hashed_p1_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23766 = _T_23243 ? bht_bank_rd_data_out_1_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24021 = _T_24020 | _T_23766; // @[Mux.scala 27:72]
  wire  _T_23246 = bht_rd_addr_hashed_p1_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23767 = _T_23246 ? bht_bank_rd_data_out_1_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24022 = _T_24021 | _T_23767; // @[Mux.scala 27:72]
  wire  _T_23249 = bht_rd_addr_hashed_p1_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23768 = _T_23249 ? bht_bank_rd_data_out_1_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24023 = _T_24022 | _T_23768; // @[Mux.scala 27:72]
  wire  _T_23252 = bht_rd_addr_hashed_p1_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23769 = _T_23252 ? bht_bank_rd_data_out_1_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24024 = _T_24023 | _T_23769; // @[Mux.scala 27:72]
  wire  _T_23255 = bht_rd_addr_hashed_p1_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23770 = _T_23255 ? bht_bank_rd_data_out_1_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24025 = _T_24024 | _T_23770; // @[Mux.scala 27:72]
  wire  _T_23258 = bht_rd_addr_hashed_p1_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23771 = _T_23258 ? bht_bank_rd_data_out_1_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24026 = _T_24025 | _T_23771; // @[Mux.scala 27:72]
  wire  _T_23261 = bht_rd_addr_hashed_p1_f == 8'h80; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23772 = _T_23261 ? bht_bank_rd_data_out_1_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24027 = _T_24026 | _T_23772; // @[Mux.scala 27:72]
  wire  _T_23264 = bht_rd_addr_hashed_p1_f == 8'h81; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23773 = _T_23264 ? bht_bank_rd_data_out_1_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24028 = _T_24027 | _T_23773; // @[Mux.scala 27:72]
  wire  _T_23267 = bht_rd_addr_hashed_p1_f == 8'h82; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23774 = _T_23267 ? bht_bank_rd_data_out_1_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24029 = _T_24028 | _T_23774; // @[Mux.scala 27:72]
  wire  _T_23270 = bht_rd_addr_hashed_p1_f == 8'h83; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23775 = _T_23270 ? bht_bank_rd_data_out_1_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24030 = _T_24029 | _T_23775; // @[Mux.scala 27:72]
  wire  _T_23273 = bht_rd_addr_hashed_p1_f == 8'h84; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23776 = _T_23273 ? bht_bank_rd_data_out_1_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24031 = _T_24030 | _T_23776; // @[Mux.scala 27:72]
  wire  _T_23276 = bht_rd_addr_hashed_p1_f == 8'h85; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23777 = _T_23276 ? bht_bank_rd_data_out_1_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24032 = _T_24031 | _T_23777; // @[Mux.scala 27:72]
  wire  _T_23279 = bht_rd_addr_hashed_p1_f == 8'h86; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23778 = _T_23279 ? bht_bank_rd_data_out_1_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24033 = _T_24032 | _T_23778; // @[Mux.scala 27:72]
  wire  _T_23282 = bht_rd_addr_hashed_p1_f == 8'h87; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23779 = _T_23282 ? bht_bank_rd_data_out_1_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24034 = _T_24033 | _T_23779; // @[Mux.scala 27:72]
  wire  _T_23285 = bht_rd_addr_hashed_p1_f == 8'h88; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23780 = _T_23285 ? bht_bank_rd_data_out_1_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24035 = _T_24034 | _T_23780; // @[Mux.scala 27:72]
  wire  _T_23288 = bht_rd_addr_hashed_p1_f == 8'h89; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23781 = _T_23288 ? bht_bank_rd_data_out_1_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24036 = _T_24035 | _T_23781; // @[Mux.scala 27:72]
  wire  _T_23291 = bht_rd_addr_hashed_p1_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23782 = _T_23291 ? bht_bank_rd_data_out_1_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24037 = _T_24036 | _T_23782; // @[Mux.scala 27:72]
  wire  _T_23294 = bht_rd_addr_hashed_p1_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23783 = _T_23294 ? bht_bank_rd_data_out_1_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24038 = _T_24037 | _T_23783; // @[Mux.scala 27:72]
  wire  _T_23297 = bht_rd_addr_hashed_p1_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23784 = _T_23297 ? bht_bank_rd_data_out_1_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24039 = _T_24038 | _T_23784; // @[Mux.scala 27:72]
  wire  _T_23300 = bht_rd_addr_hashed_p1_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23785 = _T_23300 ? bht_bank_rd_data_out_1_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24040 = _T_24039 | _T_23785; // @[Mux.scala 27:72]
  wire  _T_23303 = bht_rd_addr_hashed_p1_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23786 = _T_23303 ? bht_bank_rd_data_out_1_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24041 = _T_24040 | _T_23786; // @[Mux.scala 27:72]
  wire  _T_23306 = bht_rd_addr_hashed_p1_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23787 = _T_23306 ? bht_bank_rd_data_out_1_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24042 = _T_24041 | _T_23787; // @[Mux.scala 27:72]
  wire  _T_23309 = bht_rd_addr_hashed_p1_f == 8'h90; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23788 = _T_23309 ? bht_bank_rd_data_out_1_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24043 = _T_24042 | _T_23788; // @[Mux.scala 27:72]
  wire  _T_23312 = bht_rd_addr_hashed_p1_f == 8'h91; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23789 = _T_23312 ? bht_bank_rd_data_out_1_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24044 = _T_24043 | _T_23789; // @[Mux.scala 27:72]
  wire  _T_23315 = bht_rd_addr_hashed_p1_f == 8'h92; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23790 = _T_23315 ? bht_bank_rd_data_out_1_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24045 = _T_24044 | _T_23790; // @[Mux.scala 27:72]
  wire  _T_23318 = bht_rd_addr_hashed_p1_f == 8'h93; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23791 = _T_23318 ? bht_bank_rd_data_out_1_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24046 = _T_24045 | _T_23791; // @[Mux.scala 27:72]
  wire  _T_23321 = bht_rd_addr_hashed_p1_f == 8'h94; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23792 = _T_23321 ? bht_bank_rd_data_out_1_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24047 = _T_24046 | _T_23792; // @[Mux.scala 27:72]
  wire  _T_23324 = bht_rd_addr_hashed_p1_f == 8'h95; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23793 = _T_23324 ? bht_bank_rd_data_out_1_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24048 = _T_24047 | _T_23793; // @[Mux.scala 27:72]
  wire  _T_23327 = bht_rd_addr_hashed_p1_f == 8'h96; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23794 = _T_23327 ? bht_bank_rd_data_out_1_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24049 = _T_24048 | _T_23794; // @[Mux.scala 27:72]
  wire  _T_23330 = bht_rd_addr_hashed_p1_f == 8'h97; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23795 = _T_23330 ? bht_bank_rd_data_out_1_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24050 = _T_24049 | _T_23795; // @[Mux.scala 27:72]
  wire  _T_23333 = bht_rd_addr_hashed_p1_f == 8'h98; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23796 = _T_23333 ? bht_bank_rd_data_out_1_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24051 = _T_24050 | _T_23796; // @[Mux.scala 27:72]
  wire  _T_23336 = bht_rd_addr_hashed_p1_f == 8'h99; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23797 = _T_23336 ? bht_bank_rd_data_out_1_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24052 = _T_24051 | _T_23797; // @[Mux.scala 27:72]
  wire  _T_23339 = bht_rd_addr_hashed_p1_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23798 = _T_23339 ? bht_bank_rd_data_out_1_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24053 = _T_24052 | _T_23798; // @[Mux.scala 27:72]
  wire  _T_23342 = bht_rd_addr_hashed_p1_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23799 = _T_23342 ? bht_bank_rd_data_out_1_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24054 = _T_24053 | _T_23799; // @[Mux.scala 27:72]
  wire  _T_23345 = bht_rd_addr_hashed_p1_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23800 = _T_23345 ? bht_bank_rd_data_out_1_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24055 = _T_24054 | _T_23800; // @[Mux.scala 27:72]
  wire  _T_23348 = bht_rd_addr_hashed_p1_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23801 = _T_23348 ? bht_bank_rd_data_out_1_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24056 = _T_24055 | _T_23801; // @[Mux.scala 27:72]
  wire  _T_23351 = bht_rd_addr_hashed_p1_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23802 = _T_23351 ? bht_bank_rd_data_out_1_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24057 = _T_24056 | _T_23802; // @[Mux.scala 27:72]
  wire  _T_23354 = bht_rd_addr_hashed_p1_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23803 = _T_23354 ? bht_bank_rd_data_out_1_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24058 = _T_24057 | _T_23803; // @[Mux.scala 27:72]
  wire  _T_23357 = bht_rd_addr_hashed_p1_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23804 = _T_23357 ? bht_bank_rd_data_out_1_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24059 = _T_24058 | _T_23804; // @[Mux.scala 27:72]
  wire  _T_23360 = bht_rd_addr_hashed_p1_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23805 = _T_23360 ? bht_bank_rd_data_out_1_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24060 = _T_24059 | _T_23805; // @[Mux.scala 27:72]
  wire  _T_23363 = bht_rd_addr_hashed_p1_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23806 = _T_23363 ? bht_bank_rd_data_out_1_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24061 = _T_24060 | _T_23806; // @[Mux.scala 27:72]
  wire  _T_23366 = bht_rd_addr_hashed_p1_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23807 = _T_23366 ? bht_bank_rd_data_out_1_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24062 = _T_24061 | _T_23807; // @[Mux.scala 27:72]
  wire  _T_23369 = bht_rd_addr_hashed_p1_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23808 = _T_23369 ? bht_bank_rd_data_out_1_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24063 = _T_24062 | _T_23808; // @[Mux.scala 27:72]
  wire  _T_23372 = bht_rd_addr_hashed_p1_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23809 = _T_23372 ? bht_bank_rd_data_out_1_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24064 = _T_24063 | _T_23809; // @[Mux.scala 27:72]
  wire  _T_23375 = bht_rd_addr_hashed_p1_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23810 = _T_23375 ? bht_bank_rd_data_out_1_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24065 = _T_24064 | _T_23810; // @[Mux.scala 27:72]
  wire  _T_23378 = bht_rd_addr_hashed_p1_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23811 = _T_23378 ? bht_bank_rd_data_out_1_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24066 = _T_24065 | _T_23811; // @[Mux.scala 27:72]
  wire  _T_23381 = bht_rd_addr_hashed_p1_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23812 = _T_23381 ? bht_bank_rd_data_out_1_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24067 = _T_24066 | _T_23812; // @[Mux.scala 27:72]
  wire  _T_23384 = bht_rd_addr_hashed_p1_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23813 = _T_23384 ? bht_bank_rd_data_out_1_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24068 = _T_24067 | _T_23813; // @[Mux.scala 27:72]
  wire  _T_23387 = bht_rd_addr_hashed_p1_f == 8'haa; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23814 = _T_23387 ? bht_bank_rd_data_out_1_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24069 = _T_24068 | _T_23814; // @[Mux.scala 27:72]
  wire  _T_23390 = bht_rd_addr_hashed_p1_f == 8'hab; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23815 = _T_23390 ? bht_bank_rd_data_out_1_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24070 = _T_24069 | _T_23815; // @[Mux.scala 27:72]
  wire  _T_23393 = bht_rd_addr_hashed_p1_f == 8'hac; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23816 = _T_23393 ? bht_bank_rd_data_out_1_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24071 = _T_24070 | _T_23816; // @[Mux.scala 27:72]
  wire  _T_23396 = bht_rd_addr_hashed_p1_f == 8'had; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23817 = _T_23396 ? bht_bank_rd_data_out_1_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24072 = _T_24071 | _T_23817; // @[Mux.scala 27:72]
  wire  _T_23399 = bht_rd_addr_hashed_p1_f == 8'hae; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23818 = _T_23399 ? bht_bank_rd_data_out_1_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24073 = _T_24072 | _T_23818; // @[Mux.scala 27:72]
  wire  _T_23402 = bht_rd_addr_hashed_p1_f == 8'haf; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23819 = _T_23402 ? bht_bank_rd_data_out_1_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24074 = _T_24073 | _T_23819; // @[Mux.scala 27:72]
  wire  _T_23405 = bht_rd_addr_hashed_p1_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23820 = _T_23405 ? bht_bank_rd_data_out_1_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24075 = _T_24074 | _T_23820; // @[Mux.scala 27:72]
  wire  _T_23408 = bht_rd_addr_hashed_p1_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23821 = _T_23408 ? bht_bank_rd_data_out_1_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24076 = _T_24075 | _T_23821; // @[Mux.scala 27:72]
  wire  _T_23411 = bht_rd_addr_hashed_p1_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23822 = _T_23411 ? bht_bank_rd_data_out_1_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24077 = _T_24076 | _T_23822; // @[Mux.scala 27:72]
  wire  _T_23414 = bht_rd_addr_hashed_p1_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23823 = _T_23414 ? bht_bank_rd_data_out_1_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24078 = _T_24077 | _T_23823; // @[Mux.scala 27:72]
  wire  _T_23417 = bht_rd_addr_hashed_p1_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23824 = _T_23417 ? bht_bank_rd_data_out_1_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24079 = _T_24078 | _T_23824; // @[Mux.scala 27:72]
  wire  _T_23420 = bht_rd_addr_hashed_p1_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23825 = _T_23420 ? bht_bank_rd_data_out_1_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24080 = _T_24079 | _T_23825; // @[Mux.scala 27:72]
  wire  _T_23423 = bht_rd_addr_hashed_p1_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23826 = _T_23423 ? bht_bank_rd_data_out_1_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24081 = _T_24080 | _T_23826; // @[Mux.scala 27:72]
  wire  _T_23426 = bht_rd_addr_hashed_p1_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23827 = _T_23426 ? bht_bank_rd_data_out_1_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24082 = _T_24081 | _T_23827; // @[Mux.scala 27:72]
  wire  _T_23429 = bht_rd_addr_hashed_p1_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23828 = _T_23429 ? bht_bank_rd_data_out_1_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24083 = _T_24082 | _T_23828; // @[Mux.scala 27:72]
  wire  _T_23432 = bht_rd_addr_hashed_p1_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23829 = _T_23432 ? bht_bank_rd_data_out_1_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24084 = _T_24083 | _T_23829; // @[Mux.scala 27:72]
  wire  _T_23435 = bht_rd_addr_hashed_p1_f == 8'hba; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23830 = _T_23435 ? bht_bank_rd_data_out_1_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24085 = _T_24084 | _T_23830; // @[Mux.scala 27:72]
  wire  _T_23438 = bht_rd_addr_hashed_p1_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23831 = _T_23438 ? bht_bank_rd_data_out_1_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24086 = _T_24085 | _T_23831; // @[Mux.scala 27:72]
  wire  _T_23441 = bht_rd_addr_hashed_p1_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23832 = _T_23441 ? bht_bank_rd_data_out_1_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24087 = _T_24086 | _T_23832; // @[Mux.scala 27:72]
  wire  _T_23444 = bht_rd_addr_hashed_p1_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23833 = _T_23444 ? bht_bank_rd_data_out_1_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24088 = _T_24087 | _T_23833; // @[Mux.scala 27:72]
  wire  _T_23447 = bht_rd_addr_hashed_p1_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23834 = _T_23447 ? bht_bank_rd_data_out_1_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24089 = _T_24088 | _T_23834; // @[Mux.scala 27:72]
  wire  _T_23450 = bht_rd_addr_hashed_p1_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23835 = _T_23450 ? bht_bank_rd_data_out_1_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24090 = _T_24089 | _T_23835; // @[Mux.scala 27:72]
  wire  _T_23453 = bht_rd_addr_hashed_p1_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23836 = _T_23453 ? bht_bank_rd_data_out_1_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24091 = _T_24090 | _T_23836; // @[Mux.scala 27:72]
  wire  _T_23456 = bht_rd_addr_hashed_p1_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23837 = _T_23456 ? bht_bank_rd_data_out_1_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24092 = _T_24091 | _T_23837; // @[Mux.scala 27:72]
  wire  _T_23459 = bht_rd_addr_hashed_p1_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23838 = _T_23459 ? bht_bank_rd_data_out_1_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24093 = _T_24092 | _T_23838; // @[Mux.scala 27:72]
  wire  _T_23462 = bht_rd_addr_hashed_p1_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23839 = _T_23462 ? bht_bank_rd_data_out_1_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24094 = _T_24093 | _T_23839; // @[Mux.scala 27:72]
  wire  _T_23465 = bht_rd_addr_hashed_p1_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23840 = _T_23465 ? bht_bank_rd_data_out_1_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24095 = _T_24094 | _T_23840; // @[Mux.scala 27:72]
  wire  _T_23468 = bht_rd_addr_hashed_p1_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23841 = _T_23468 ? bht_bank_rd_data_out_1_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24096 = _T_24095 | _T_23841; // @[Mux.scala 27:72]
  wire  _T_23471 = bht_rd_addr_hashed_p1_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23842 = _T_23471 ? bht_bank_rd_data_out_1_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24097 = _T_24096 | _T_23842; // @[Mux.scala 27:72]
  wire  _T_23474 = bht_rd_addr_hashed_p1_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23843 = _T_23474 ? bht_bank_rd_data_out_1_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24098 = _T_24097 | _T_23843; // @[Mux.scala 27:72]
  wire  _T_23477 = bht_rd_addr_hashed_p1_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23844 = _T_23477 ? bht_bank_rd_data_out_1_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24099 = _T_24098 | _T_23844; // @[Mux.scala 27:72]
  wire  _T_23480 = bht_rd_addr_hashed_p1_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23845 = _T_23480 ? bht_bank_rd_data_out_1_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24100 = _T_24099 | _T_23845; // @[Mux.scala 27:72]
  wire  _T_23483 = bht_rd_addr_hashed_p1_f == 8'hca; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23846 = _T_23483 ? bht_bank_rd_data_out_1_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24101 = _T_24100 | _T_23846; // @[Mux.scala 27:72]
  wire  _T_23486 = bht_rd_addr_hashed_p1_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23847 = _T_23486 ? bht_bank_rd_data_out_1_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24102 = _T_24101 | _T_23847; // @[Mux.scala 27:72]
  wire  _T_23489 = bht_rd_addr_hashed_p1_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23848 = _T_23489 ? bht_bank_rd_data_out_1_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24103 = _T_24102 | _T_23848; // @[Mux.scala 27:72]
  wire  _T_23492 = bht_rd_addr_hashed_p1_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23849 = _T_23492 ? bht_bank_rd_data_out_1_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24104 = _T_24103 | _T_23849; // @[Mux.scala 27:72]
  wire  _T_23495 = bht_rd_addr_hashed_p1_f == 8'hce; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23850 = _T_23495 ? bht_bank_rd_data_out_1_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24105 = _T_24104 | _T_23850; // @[Mux.scala 27:72]
  wire  _T_23498 = bht_rd_addr_hashed_p1_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23851 = _T_23498 ? bht_bank_rd_data_out_1_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24106 = _T_24105 | _T_23851; // @[Mux.scala 27:72]
  wire  _T_23501 = bht_rd_addr_hashed_p1_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23852 = _T_23501 ? bht_bank_rd_data_out_1_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24107 = _T_24106 | _T_23852; // @[Mux.scala 27:72]
  wire  _T_23504 = bht_rd_addr_hashed_p1_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23853 = _T_23504 ? bht_bank_rd_data_out_1_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24108 = _T_24107 | _T_23853; // @[Mux.scala 27:72]
  wire  _T_23507 = bht_rd_addr_hashed_p1_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23854 = _T_23507 ? bht_bank_rd_data_out_1_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24109 = _T_24108 | _T_23854; // @[Mux.scala 27:72]
  wire  _T_23510 = bht_rd_addr_hashed_p1_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23855 = _T_23510 ? bht_bank_rd_data_out_1_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24110 = _T_24109 | _T_23855; // @[Mux.scala 27:72]
  wire  _T_23513 = bht_rd_addr_hashed_p1_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23856 = _T_23513 ? bht_bank_rd_data_out_1_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24111 = _T_24110 | _T_23856; // @[Mux.scala 27:72]
  wire  _T_23516 = bht_rd_addr_hashed_p1_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23857 = _T_23516 ? bht_bank_rd_data_out_1_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24112 = _T_24111 | _T_23857; // @[Mux.scala 27:72]
  wire  _T_23519 = bht_rd_addr_hashed_p1_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23858 = _T_23519 ? bht_bank_rd_data_out_1_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24113 = _T_24112 | _T_23858; // @[Mux.scala 27:72]
  wire  _T_23522 = bht_rd_addr_hashed_p1_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23859 = _T_23522 ? bht_bank_rd_data_out_1_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24114 = _T_24113 | _T_23859; // @[Mux.scala 27:72]
  wire  _T_23525 = bht_rd_addr_hashed_p1_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23860 = _T_23525 ? bht_bank_rd_data_out_1_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24115 = _T_24114 | _T_23860; // @[Mux.scala 27:72]
  wire  _T_23528 = bht_rd_addr_hashed_p1_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23861 = _T_23528 ? bht_bank_rd_data_out_1_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24116 = _T_24115 | _T_23861; // @[Mux.scala 27:72]
  wire  _T_23531 = bht_rd_addr_hashed_p1_f == 8'hda; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23862 = _T_23531 ? bht_bank_rd_data_out_1_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24117 = _T_24116 | _T_23862; // @[Mux.scala 27:72]
  wire  _T_23534 = bht_rd_addr_hashed_p1_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23863 = _T_23534 ? bht_bank_rd_data_out_1_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24118 = _T_24117 | _T_23863; // @[Mux.scala 27:72]
  wire  _T_23537 = bht_rd_addr_hashed_p1_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23864 = _T_23537 ? bht_bank_rd_data_out_1_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24119 = _T_24118 | _T_23864; // @[Mux.scala 27:72]
  wire  _T_23540 = bht_rd_addr_hashed_p1_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23865 = _T_23540 ? bht_bank_rd_data_out_1_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24120 = _T_24119 | _T_23865; // @[Mux.scala 27:72]
  wire  _T_23543 = bht_rd_addr_hashed_p1_f == 8'hde; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23866 = _T_23543 ? bht_bank_rd_data_out_1_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24121 = _T_24120 | _T_23866; // @[Mux.scala 27:72]
  wire  _T_23546 = bht_rd_addr_hashed_p1_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23867 = _T_23546 ? bht_bank_rd_data_out_1_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24122 = _T_24121 | _T_23867; // @[Mux.scala 27:72]
  wire  _T_23549 = bht_rd_addr_hashed_p1_f == 8'he0; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23868 = _T_23549 ? bht_bank_rd_data_out_1_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24123 = _T_24122 | _T_23868; // @[Mux.scala 27:72]
  wire  _T_23552 = bht_rd_addr_hashed_p1_f == 8'he1; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23869 = _T_23552 ? bht_bank_rd_data_out_1_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24124 = _T_24123 | _T_23869; // @[Mux.scala 27:72]
  wire  _T_23555 = bht_rd_addr_hashed_p1_f == 8'he2; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23870 = _T_23555 ? bht_bank_rd_data_out_1_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24125 = _T_24124 | _T_23870; // @[Mux.scala 27:72]
  wire  _T_23558 = bht_rd_addr_hashed_p1_f == 8'he3; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23871 = _T_23558 ? bht_bank_rd_data_out_1_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24126 = _T_24125 | _T_23871; // @[Mux.scala 27:72]
  wire  _T_23561 = bht_rd_addr_hashed_p1_f == 8'he4; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23872 = _T_23561 ? bht_bank_rd_data_out_1_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24127 = _T_24126 | _T_23872; // @[Mux.scala 27:72]
  wire  _T_23564 = bht_rd_addr_hashed_p1_f == 8'he5; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23873 = _T_23564 ? bht_bank_rd_data_out_1_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24128 = _T_24127 | _T_23873; // @[Mux.scala 27:72]
  wire  _T_23567 = bht_rd_addr_hashed_p1_f == 8'he6; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23874 = _T_23567 ? bht_bank_rd_data_out_1_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24129 = _T_24128 | _T_23874; // @[Mux.scala 27:72]
  wire  _T_23570 = bht_rd_addr_hashed_p1_f == 8'he7; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23875 = _T_23570 ? bht_bank_rd_data_out_1_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24130 = _T_24129 | _T_23875; // @[Mux.scala 27:72]
  wire  _T_23573 = bht_rd_addr_hashed_p1_f == 8'he8; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23876 = _T_23573 ? bht_bank_rd_data_out_1_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24131 = _T_24130 | _T_23876; // @[Mux.scala 27:72]
  wire  _T_23576 = bht_rd_addr_hashed_p1_f == 8'he9; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23877 = _T_23576 ? bht_bank_rd_data_out_1_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24132 = _T_24131 | _T_23877; // @[Mux.scala 27:72]
  wire  _T_23579 = bht_rd_addr_hashed_p1_f == 8'hea; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23878 = _T_23579 ? bht_bank_rd_data_out_1_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24133 = _T_24132 | _T_23878; // @[Mux.scala 27:72]
  wire  _T_23582 = bht_rd_addr_hashed_p1_f == 8'heb; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23879 = _T_23582 ? bht_bank_rd_data_out_1_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24134 = _T_24133 | _T_23879; // @[Mux.scala 27:72]
  wire  _T_23585 = bht_rd_addr_hashed_p1_f == 8'hec; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23880 = _T_23585 ? bht_bank_rd_data_out_1_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24135 = _T_24134 | _T_23880; // @[Mux.scala 27:72]
  wire  _T_23588 = bht_rd_addr_hashed_p1_f == 8'hed; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23881 = _T_23588 ? bht_bank_rd_data_out_1_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24136 = _T_24135 | _T_23881; // @[Mux.scala 27:72]
  wire  _T_23591 = bht_rd_addr_hashed_p1_f == 8'hee; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23882 = _T_23591 ? bht_bank_rd_data_out_1_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24137 = _T_24136 | _T_23882; // @[Mux.scala 27:72]
  wire  _T_23594 = bht_rd_addr_hashed_p1_f == 8'hef; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23883 = _T_23594 ? bht_bank_rd_data_out_1_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24138 = _T_24137 | _T_23883; // @[Mux.scala 27:72]
  wire  _T_23597 = bht_rd_addr_hashed_p1_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23884 = _T_23597 ? bht_bank_rd_data_out_1_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24139 = _T_24138 | _T_23884; // @[Mux.scala 27:72]
  wire  _T_23600 = bht_rd_addr_hashed_p1_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23885 = _T_23600 ? bht_bank_rd_data_out_1_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24140 = _T_24139 | _T_23885; // @[Mux.scala 27:72]
  wire  _T_23603 = bht_rd_addr_hashed_p1_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23886 = _T_23603 ? bht_bank_rd_data_out_1_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24141 = _T_24140 | _T_23886; // @[Mux.scala 27:72]
  wire  _T_23606 = bht_rd_addr_hashed_p1_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23887 = _T_23606 ? bht_bank_rd_data_out_1_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24142 = _T_24141 | _T_23887; // @[Mux.scala 27:72]
  wire  _T_23609 = bht_rd_addr_hashed_p1_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23888 = _T_23609 ? bht_bank_rd_data_out_1_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24143 = _T_24142 | _T_23888; // @[Mux.scala 27:72]
  wire  _T_23612 = bht_rd_addr_hashed_p1_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23889 = _T_23612 ? bht_bank_rd_data_out_1_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24144 = _T_24143 | _T_23889; // @[Mux.scala 27:72]
  wire  _T_23615 = bht_rd_addr_hashed_p1_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23890 = _T_23615 ? bht_bank_rd_data_out_1_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24145 = _T_24144 | _T_23890; // @[Mux.scala 27:72]
  wire  _T_23618 = bht_rd_addr_hashed_p1_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23891 = _T_23618 ? bht_bank_rd_data_out_1_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24146 = _T_24145 | _T_23891; // @[Mux.scala 27:72]
  wire  _T_23621 = bht_rd_addr_hashed_p1_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23892 = _T_23621 ? bht_bank_rd_data_out_1_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24147 = _T_24146 | _T_23892; // @[Mux.scala 27:72]
  wire  _T_23624 = bht_rd_addr_hashed_p1_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23893 = _T_23624 ? bht_bank_rd_data_out_1_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24148 = _T_24147 | _T_23893; // @[Mux.scala 27:72]
  wire  _T_23627 = bht_rd_addr_hashed_p1_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23894 = _T_23627 ? bht_bank_rd_data_out_1_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24149 = _T_24148 | _T_23894; // @[Mux.scala 27:72]
  wire  _T_23630 = bht_rd_addr_hashed_p1_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23895 = _T_23630 ? bht_bank_rd_data_out_1_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24150 = _T_24149 | _T_23895; // @[Mux.scala 27:72]
  wire  _T_23633 = bht_rd_addr_hashed_p1_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23896 = _T_23633 ? bht_bank_rd_data_out_1_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24151 = _T_24150 | _T_23896; // @[Mux.scala 27:72]
  wire  _T_23636 = bht_rd_addr_hashed_p1_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23897 = _T_23636 ? bht_bank_rd_data_out_1_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24152 = _T_24151 | _T_23897; // @[Mux.scala 27:72]
  wire  _T_23639 = bht_rd_addr_hashed_p1_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23898 = _T_23639 ? bht_bank_rd_data_out_1_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24153 = _T_24152 | _T_23898; // @[Mux.scala 27:72]
  wire  _T_23642 = bht_rd_addr_hashed_p1_f == 8'hff; // @[el2_ifu_bp_ctl.scala 397:112]
  wire [1:0] _T_23899 = _T_23642 ? bht_bank_rd_data_out_1_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_p1_f = _T_24153 | _T_23899; // @[Mux.scala 27:72]
  wire [1:0] _T_259 = io_ifc_fetch_addr_f[0] ? bht_bank0_rd_data_p1_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank1_rd_data_f = _T_258 | _T_259; // @[Mux.scala 27:72]
  wire  _T_263 = bht_force_taken_f[1] | bht_vbank1_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 250:42]
  wire [1:0] wayhit_f = tag_match_way0_expanded_f | tag_match_way1_expanded_f; // @[el2_ifu_bp_ctl.scala 160:44]
  wire [1:0] _T_158 = _T_143 ? wayhit_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] wayhit_p1_f = tag_match_way0_expanded_p1_f | tag_match_way1_expanded_p1_f; // @[el2_ifu_bp_ctl.scala 162:50]
  wire [1:0] _T_157 = {wayhit_p1_f[0],wayhit_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_159 = io_ifc_fetch_addr_f[0] ? _T_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_160 = _T_158 | _T_159; // @[Mux.scala 27:72]
  wire  eoc_near = &io_ifc_fetch_addr_f[4:2]; // @[el2_ifu_bp_ctl.scala 219:64]
  wire  _T_217 = ~eoc_near; // @[el2_ifu_bp_ctl.scala 221:15]
  wire  _T_219 = |io_ifc_fetch_addr_f[1:0]; // @[el2_ifu_bp_ctl.scala 221:57]
  wire  _T_220 = ~_T_219; // @[el2_ifu_bp_ctl.scala 221:28]
  wire  eoc_mask = _T_217 | _T_220; // @[el2_ifu_bp_ctl.scala 221:25]
  wire [1:0] _T_162 = {eoc_mask,1'h1}; // @[Cat.scala 29:58]
  wire [1:0] vwayhit_f = _T_160 & _T_162; // @[el2_ifu_bp_ctl.scala 189:71]
  wire  _T_265 = _T_263 & vwayhit_f[1]; // @[el2_ifu_bp_ctl.scala 250:69]
  reg [1:0] bht_bank_rd_data_out_0_0; // @[Reg.scala 27:20]
  wire [1:0] _T_21084 = _T_21597 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_1; // @[Reg.scala 27:20]
  wire [1:0] _T_21085 = _T_21600 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21340 = _T_21084 | _T_21085; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_2; // @[Reg.scala 27:20]
  wire [1:0] _T_21086 = _T_21603 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21341 = _T_21340 | _T_21086; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_3; // @[Reg.scala 27:20]
  wire [1:0] _T_21087 = _T_21606 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21342 = _T_21341 | _T_21087; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_4; // @[Reg.scala 27:20]
  wire [1:0] _T_21088 = _T_21609 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21343 = _T_21342 | _T_21088; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_5; // @[Reg.scala 27:20]
  wire [1:0] _T_21089 = _T_21612 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21344 = _T_21343 | _T_21089; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_6; // @[Reg.scala 27:20]
  wire [1:0] _T_21090 = _T_21615 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21345 = _T_21344 | _T_21090; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_7; // @[Reg.scala 27:20]
  wire [1:0] _T_21091 = _T_21618 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21346 = _T_21345 | _T_21091; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_8; // @[Reg.scala 27:20]
  wire [1:0] _T_21092 = _T_21621 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21347 = _T_21346 | _T_21092; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_9; // @[Reg.scala 27:20]
  wire [1:0] _T_21093 = _T_21624 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21348 = _T_21347 | _T_21093; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_10; // @[Reg.scala 27:20]
  wire [1:0] _T_21094 = _T_21627 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21349 = _T_21348 | _T_21094; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_11; // @[Reg.scala 27:20]
  wire [1:0] _T_21095 = _T_21630 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21350 = _T_21349 | _T_21095; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_12; // @[Reg.scala 27:20]
  wire [1:0] _T_21096 = _T_21633 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21351 = _T_21350 | _T_21096; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_13; // @[Reg.scala 27:20]
  wire [1:0] _T_21097 = _T_21636 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21352 = _T_21351 | _T_21097; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_14; // @[Reg.scala 27:20]
  wire [1:0] _T_21098 = _T_21639 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21353 = _T_21352 | _T_21098; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_15; // @[Reg.scala 27:20]
  wire [1:0] _T_21099 = _T_21642 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21354 = _T_21353 | _T_21099; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_16; // @[Reg.scala 27:20]
  wire [1:0] _T_21100 = _T_21645 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21355 = _T_21354 | _T_21100; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_17; // @[Reg.scala 27:20]
  wire [1:0] _T_21101 = _T_21648 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21356 = _T_21355 | _T_21101; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_18; // @[Reg.scala 27:20]
  wire [1:0] _T_21102 = _T_21651 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21357 = _T_21356 | _T_21102; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_19; // @[Reg.scala 27:20]
  wire [1:0] _T_21103 = _T_21654 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21358 = _T_21357 | _T_21103; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_20; // @[Reg.scala 27:20]
  wire [1:0] _T_21104 = _T_21657 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21359 = _T_21358 | _T_21104; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_21; // @[Reg.scala 27:20]
  wire [1:0] _T_21105 = _T_21660 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21360 = _T_21359 | _T_21105; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_22; // @[Reg.scala 27:20]
  wire [1:0] _T_21106 = _T_21663 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21361 = _T_21360 | _T_21106; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_23; // @[Reg.scala 27:20]
  wire [1:0] _T_21107 = _T_21666 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21362 = _T_21361 | _T_21107; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_24; // @[Reg.scala 27:20]
  wire [1:0] _T_21108 = _T_21669 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21363 = _T_21362 | _T_21108; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_25; // @[Reg.scala 27:20]
  wire [1:0] _T_21109 = _T_21672 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21364 = _T_21363 | _T_21109; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_26; // @[Reg.scala 27:20]
  wire [1:0] _T_21110 = _T_21675 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21365 = _T_21364 | _T_21110; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_27; // @[Reg.scala 27:20]
  wire [1:0] _T_21111 = _T_21678 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21366 = _T_21365 | _T_21111; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_28; // @[Reg.scala 27:20]
  wire [1:0] _T_21112 = _T_21681 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21367 = _T_21366 | _T_21112; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_29; // @[Reg.scala 27:20]
  wire [1:0] _T_21113 = _T_21684 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21368 = _T_21367 | _T_21113; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_30; // @[Reg.scala 27:20]
  wire [1:0] _T_21114 = _T_21687 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21369 = _T_21368 | _T_21114; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_31; // @[Reg.scala 27:20]
  wire [1:0] _T_21115 = _T_21690 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21370 = _T_21369 | _T_21115; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_32; // @[Reg.scala 27:20]
  wire [1:0] _T_21116 = _T_21693 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21371 = _T_21370 | _T_21116; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_33; // @[Reg.scala 27:20]
  wire [1:0] _T_21117 = _T_21696 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21372 = _T_21371 | _T_21117; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_34; // @[Reg.scala 27:20]
  wire [1:0] _T_21118 = _T_21699 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21373 = _T_21372 | _T_21118; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_35; // @[Reg.scala 27:20]
  wire [1:0] _T_21119 = _T_21702 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21374 = _T_21373 | _T_21119; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_36; // @[Reg.scala 27:20]
  wire [1:0] _T_21120 = _T_21705 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21375 = _T_21374 | _T_21120; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_37; // @[Reg.scala 27:20]
  wire [1:0] _T_21121 = _T_21708 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21376 = _T_21375 | _T_21121; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_38; // @[Reg.scala 27:20]
  wire [1:0] _T_21122 = _T_21711 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21377 = _T_21376 | _T_21122; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_39; // @[Reg.scala 27:20]
  wire [1:0] _T_21123 = _T_21714 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21378 = _T_21377 | _T_21123; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_40; // @[Reg.scala 27:20]
  wire [1:0] _T_21124 = _T_21717 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21379 = _T_21378 | _T_21124; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_41; // @[Reg.scala 27:20]
  wire [1:0] _T_21125 = _T_21720 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21380 = _T_21379 | _T_21125; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_42; // @[Reg.scala 27:20]
  wire [1:0] _T_21126 = _T_21723 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21381 = _T_21380 | _T_21126; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_43; // @[Reg.scala 27:20]
  wire [1:0] _T_21127 = _T_21726 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21382 = _T_21381 | _T_21127; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_44; // @[Reg.scala 27:20]
  wire [1:0] _T_21128 = _T_21729 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21383 = _T_21382 | _T_21128; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_45; // @[Reg.scala 27:20]
  wire [1:0] _T_21129 = _T_21732 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21384 = _T_21383 | _T_21129; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_46; // @[Reg.scala 27:20]
  wire [1:0] _T_21130 = _T_21735 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21385 = _T_21384 | _T_21130; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_47; // @[Reg.scala 27:20]
  wire [1:0] _T_21131 = _T_21738 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21386 = _T_21385 | _T_21131; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_48; // @[Reg.scala 27:20]
  wire [1:0] _T_21132 = _T_21741 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21387 = _T_21386 | _T_21132; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_49; // @[Reg.scala 27:20]
  wire [1:0] _T_21133 = _T_21744 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21388 = _T_21387 | _T_21133; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_50; // @[Reg.scala 27:20]
  wire [1:0] _T_21134 = _T_21747 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21389 = _T_21388 | _T_21134; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_51; // @[Reg.scala 27:20]
  wire [1:0] _T_21135 = _T_21750 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21390 = _T_21389 | _T_21135; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_52; // @[Reg.scala 27:20]
  wire [1:0] _T_21136 = _T_21753 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21391 = _T_21390 | _T_21136; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_53; // @[Reg.scala 27:20]
  wire [1:0] _T_21137 = _T_21756 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21392 = _T_21391 | _T_21137; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_54; // @[Reg.scala 27:20]
  wire [1:0] _T_21138 = _T_21759 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21393 = _T_21392 | _T_21138; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_55; // @[Reg.scala 27:20]
  wire [1:0] _T_21139 = _T_21762 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21394 = _T_21393 | _T_21139; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_56; // @[Reg.scala 27:20]
  wire [1:0] _T_21140 = _T_21765 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21395 = _T_21394 | _T_21140; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_57; // @[Reg.scala 27:20]
  wire [1:0] _T_21141 = _T_21768 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21396 = _T_21395 | _T_21141; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_58; // @[Reg.scala 27:20]
  wire [1:0] _T_21142 = _T_21771 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21397 = _T_21396 | _T_21142; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_59; // @[Reg.scala 27:20]
  wire [1:0] _T_21143 = _T_21774 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21398 = _T_21397 | _T_21143; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_60; // @[Reg.scala 27:20]
  wire [1:0] _T_21144 = _T_21777 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21399 = _T_21398 | _T_21144; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_61; // @[Reg.scala 27:20]
  wire [1:0] _T_21145 = _T_21780 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21400 = _T_21399 | _T_21145; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_62; // @[Reg.scala 27:20]
  wire [1:0] _T_21146 = _T_21783 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21401 = _T_21400 | _T_21146; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_63; // @[Reg.scala 27:20]
  wire [1:0] _T_21147 = _T_21786 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21402 = _T_21401 | _T_21147; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_64; // @[Reg.scala 27:20]
  wire [1:0] _T_21148 = _T_21789 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21403 = _T_21402 | _T_21148; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_65; // @[Reg.scala 27:20]
  wire [1:0] _T_21149 = _T_21792 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21404 = _T_21403 | _T_21149; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_66; // @[Reg.scala 27:20]
  wire [1:0] _T_21150 = _T_21795 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21405 = _T_21404 | _T_21150; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_67; // @[Reg.scala 27:20]
  wire [1:0] _T_21151 = _T_21798 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21406 = _T_21405 | _T_21151; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_68; // @[Reg.scala 27:20]
  wire [1:0] _T_21152 = _T_21801 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21407 = _T_21406 | _T_21152; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_69; // @[Reg.scala 27:20]
  wire [1:0] _T_21153 = _T_21804 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21408 = _T_21407 | _T_21153; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_70; // @[Reg.scala 27:20]
  wire [1:0] _T_21154 = _T_21807 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21409 = _T_21408 | _T_21154; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_71; // @[Reg.scala 27:20]
  wire [1:0] _T_21155 = _T_21810 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21410 = _T_21409 | _T_21155; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_72; // @[Reg.scala 27:20]
  wire [1:0] _T_21156 = _T_21813 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21411 = _T_21410 | _T_21156; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_73; // @[Reg.scala 27:20]
  wire [1:0] _T_21157 = _T_21816 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21412 = _T_21411 | _T_21157; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_74; // @[Reg.scala 27:20]
  wire [1:0] _T_21158 = _T_21819 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21413 = _T_21412 | _T_21158; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_75; // @[Reg.scala 27:20]
  wire [1:0] _T_21159 = _T_21822 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21414 = _T_21413 | _T_21159; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_76; // @[Reg.scala 27:20]
  wire [1:0] _T_21160 = _T_21825 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21415 = _T_21414 | _T_21160; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_77; // @[Reg.scala 27:20]
  wire [1:0] _T_21161 = _T_21828 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21416 = _T_21415 | _T_21161; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_78; // @[Reg.scala 27:20]
  wire [1:0] _T_21162 = _T_21831 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21417 = _T_21416 | _T_21162; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_79; // @[Reg.scala 27:20]
  wire [1:0] _T_21163 = _T_21834 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21418 = _T_21417 | _T_21163; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_80; // @[Reg.scala 27:20]
  wire [1:0] _T_21164 = _T_21837 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21419 = _T_21418 | _T_21164; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_81; // @[Reg.scala 27:20]
  wire [1:0] _T_21165 = _T_21840 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21420 = _T_21419 | _T_21165; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_82; // @[Reg.scala 27:20]
  wire [1:0] _T_21166 = _T_21843 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21421 = _T_21420 | _T_21166; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_83; // @[Reg.scala 27:20]
  wire [1:0] _T_21167 = _T_21846 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21422 = _T_21421 | _T_21167; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_84; // @[Reg.scala 27:20]
  wire [1:0] _T_21168 = _T_21849 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21423 = _T_21422 | _T_21168; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_85; // @[Reg.scala 27:20]
  wire [1:0] _T_21169 = _T_21852 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21424 = _T_21423 | _T_21169; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_86; // @[Reg.scala 27:20]
  wire [1:0] _T_21170 = _T_21855 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21425 = _T_21424 | _T_21170; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_87; // @[Reg.scala 27:20]
  wire [1:0] _T_21171 = _T_21858 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21426 = _T_21425 | _T_21171; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_88; // @[Reg.scala 27:20]
  wire [1:0] _T_21172 = _T_21861 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21427 = _T_21426 | _T_21172; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_89; // @[Reg.scala 27:20]
  wire [1:0] _T_21173 = _T_21864 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21428 = _T_21427 | _T_21173; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_90; // @[Reg.scala 27:20]
  wire [1:0] _T_21174 = _T_21867 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21429 = _T_21428 | _T_21174; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_91; // @[Reg.scala 27:20]
  wire [1:0] _T_21175 = _T_21870 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21430 = _T_21429 | _T_21175; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_92; // @[Reg.scala 27:20]
  wire [1:0] _T_21176 = _T_21873 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21431 = _T_21430 | _T_21176; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_93; // @[Reg.scala 27:20]
  wire [1:0] _T_21177 = _T_21876 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21432 = _T_21431 | _T_21177; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_94; // @[Reg.scala 27:20]
  wire [1:0] _T_21178 = _T_21879 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21433 = _T_21432 | _T_21178; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_95; // @[Reg.scala 27:20]
  wire [1:0] _T_21179 = _T_21882 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21434 = _T_21433 | _T_21179; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_96; // @[Reg.scala 27:20]
  wire [1:0] _T_21180 = _T_21885 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21435 = _T_21434 | _T_21180; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_97; // @[Reg.scala 27:20]
  wire [1:0] _T_21181 = _T_21888 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21436 = _T_21435 | _T_21181; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_98; // @[Reg.scala 27:20]
  wire [1:0] _T_21182 = _T_21891 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21437 = _T_21436 | _T_21182; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_99; // @[Reg.scala 27:20]
  wire [1:0] _T_21183 = _T_21894 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21438 = _T_21437 | _T_21183; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_100; // @[Reg.scala 27:20]
  wire [1:0] _T_21184 = _T_21897 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21439 = _T_21438 | _T_21184; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_101; // @[Reg.scala 27:20]
  wire [1:0] _T_21185 = _T_21900 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21440 = _T_21439 | _T_21185; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_102; // @[Reg.scala 27:20]
  wire [1:0] _T_21186 = _T_21903 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21441 = _T_21440 | _T_21186; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_103; // @[Reg.scala 27:20]
  wire [1:0] _T_21187 = _T_21906 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21442 = _T_21441 | _T_21187; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_104; // @[Reg.scala 27:20]
  wire [1:0] _T_21188 = _T_21909 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21443 = _T_21442 | _T_21188; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_105; // @[Reg.scala 27:20]
  wire [1:0] _T_21189 = _T_21912 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21444 = _T_21443 | _T_21189; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_106; // @[Reg.scala 27:20]
  wire [1:0] _T_21190 = _T_21915 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21445 = _T_21444 | _T_21190; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_107; // @[Reg.scala 27:20]
  wire [1:0] _T_21191 = _T_21918 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21446 = _T_21445 | _T_21191; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_108; // @[Reg.scala 27:20]
  wire [1:0] _T_21192 = _T_21921 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21447 = _T_21446 | _T_21192; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_109; // @[Reg.scala 27:20]
  wire [1:0] _T_21193 = _T_21924 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21448 = _T_21447 | _T_21193; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_110; // @[Reg.scala 27:20]
  wire [1:0] _T_21194 = _T_21927 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21449 = _T_21448 | _T_21194; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_111; // @[Reg.scala 27:20]
  wire [1:0] _T_21195 = _T_21930 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21450 = _T_21449 | _T_21195; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_112; // @[Reg.scala 27:20]
  wire [1:0] _T_21196 = _T_21933 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21451 = _T_21450 | _T_21196; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_113; // @[Reg.scala 27:20]
  wire [1:0] _T_21197 = _T_21936 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21452 = _T_21451 | _T_21197; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_114; // @[Reg.scala 27:20]
  wire [1:0] _T_21198 = _T_21939 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21453 = _T_21452 | _T_21198; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_115; // @[Reg.scala 27:20]
  wire [1:0] _T_21199 = _T_21942 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21454 = _T_21453 | _T_21199; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_116; // @[Reg.scala 27:20]
  wire [1:0] _T_21200 = _T_21945 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21455 = _T_21454 | _T_21200; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_117; // @[Reg.scala 27:20]
  wire [1:0] _T_21201 = _T_21948 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21456 = _T_21455 | _T_21201; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_118; // @[Reg.scala 27:20]
  wire [1:0] _T_21202 = _T_21951 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21457 = _T_21456 | _T_21202; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_119; // @[Reg.scala 27:20]
  wire [1:0] _T_21203 = _T_21954 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21458 = _T_21457 | _T_21203; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_120; // @[Reg.scala 27:20]
  wire [1:0] _T_21204 = _T_21957 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21459 = _T_21458 | _T_21204; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_121; // @[Reg.scala 27:20]
  wire [1:0] _T_21205 = _T_21960 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21460 = _T_21459 | _T_21205; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_122; // @[Reg.scala 27:20]
  wire [1:0] _T_21206 = _T_21963 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21461 = _T_21460 | _T_21206; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_123; // @[Reg.scala 27:20]
  wire [1:0] _T_21207 = _T_21966 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21462 = _T_21461 | _T_21207; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_124; // @[Reg.scala 27:20]
  wire [1:0] _T_21208 = _T_21969 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21463 = _T_21462 | _T_21208; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_125; // @[Reg.scala 27:20]
  wire [1:0] _T_21209 = _T_21972 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21464 = _T_21463 | _T_21209; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_126; // @[Reg.scala 27:20]
  wire [1:0] _T_21210 = _T_21975 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21465 = _T_21464 | _T_21210; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_127; // @[Reg.scala 27:20]
  wire [1:0] _T_21211 = _T_21978 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21466 = _T_21465 | _T_21211; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_128; // @[Reg.scala 27:20]
  wire [1:0] _T_21212 = _T_21981 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21467 = _T_21466 | _T_21212; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_129; // @[Reg.scala 27:20]
  wire [1:0] _T_21213 = _T_21984 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21468 = _T_21467 | _T_21213; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_130; // @[Reg.scala 27:20]
  wire [1:0] _T_21214 = _T_21987 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21469 = _T_21468 | _T_21214; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_131; // @[Reg.scala 27:20]
  wire [1:0] _T_21215 = _T_21990 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21470 = _T_21469 | _T_21215; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_132; // @[Reg.scala 27:20]
  wire [1:0] _T_21216 = _T_21993 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21471 = _T_21470 | _T_21216; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_133; // @[Reg.scala 27:20]
  wire [1:0] _T_21217 = _T_21996 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21472 = _T_21471 | _T_21217; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_134; // @[Reg.scala 27:20]
  wire [1:0] _T_21218 = _T_21999 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21473 = _T_21472 | _T_21218; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_135; // @[Reg.scala 27:20]
  wire [1:0] _T_21219 = _T_22002 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21474 = _T_21473 | _T_21219; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_136; // @[Reg.scala 27:20]
  wire [1:0] _T_21220 = _T_22005 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21475 = _T_21474 | _T_21220; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_137; // @[Reg.scala 27:20]
  wire [1:0] _T_21221 = _T_22008 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21476 = _T_21475 | _T_21221; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_138; // @[Reg.scala 27:20]
  wire [1:0] _T_21222 = _T_22011 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21477 = _T_21476 | _T_21222; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_139; // @[Reg.scala 27:20]
  wire [1:0] _T_21223 = _T_22014 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21478 = _T_21477 | _T_21223; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_140; // @[Reg.scala 27:20]
  wire [1:0] _T_21224 = _T_22017 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21479 = _T_21478 | _T_21224; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_141; // @[Reg.scala 27:20]
  wire [1:0] _T_21225 = _T_22020 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21480 = _T_21479 | _T_21225; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_142; // @[Reg.scala 27:20]
  wire [1:0] _T_21226 = _T_22023 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21481 = _T_21480 | _T_21226; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_143; // @[Reg.scala 27:20]
  wire [1:0] _T_21227 = _T_22026 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21482 = _T_21481 | _T_21227; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_144; // @[Reg.scala 27:20]
  wire [1:0] _T_21228 = _T_22029 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21483 = _T_21482 | _T_21228; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_145; // @[Reg.scala 27:20]
  wire [1:0] _T_21229 = _T_22032 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21484 = _T_21483 | _T_21229; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_146; // @[Reg.scala 27:20]
  wire [1:0] _T_21230 = _T_22035 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21485 = _T_21484 | _T_21230; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_147; // @[Reg.scala 27:20]
  wire [1:0] _T_21231 = _T_22038 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21486 = _T_21485 | _T_21231; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_148; // @[Reg.scala 27:20]
  wire [1:0] _T_21232 = _T_22041 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21487 = _T_21486 | _T_21232; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_149; // @[Reg.scala 27:20]
  wire [1:0] _T_21233 = _T_22044 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21488 = _T_21487 | _T_21233; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_150; // @[Reg.scala 27:20]
  wire [1:0] _T_21234 = _T_22047 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21489 = _T_21488 | _T_21234; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_151; // @[Reg.scala 27:20]
  wire [1:0] _T_21235 = _T_22050 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21490 = _T_21489 | _T_21235; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_152; // @[Reg.scala 27:20]
  wire [1:0] _T_21236 = _T_22053 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21491 = _T_21490 | _T_21236; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_153; // @[Reg.scala 27:20]
  wire [1:0] _T_21237 = _T_22056 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21492 = _T_21491 | _T_21237; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_154; // @[Reg.scala 27:20]
  wire [1:0] _T_21238 = _T_22059 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21493 = _T_21492 | _T_21238; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_155; // @[Reg.scala 27:20]
  wire [1:0] _T_21239 = _T_22062 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21494 = _T_21493 | _T_21239; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_156; // @[Reg.scala 27:20]
  wire [1:0] _T_21240 = _T_22065 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21495 = _T_21494 | _T_21240; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_157; // @[Reg.scala 27:20]
  wire [1:0] _T_21241 = _T_22068 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21496 = _T_21495 | _T_21241; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_158; // @[Reg.scala 27:20]
  wire [1:0] _T_21242 = _T_22071 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21497 = _T_21496 | _T_21242; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_159; // @[Reg.scala 27:20]
  wire [1:0] _T_21243 = _T_22074 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21498 = _T_21497 | _T_21243; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_160; // @[Reg.scala 27:20]
  wire [1:0] _T_21244 = _T_22077 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21499 = _T_21498 | _T_21244; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_161; // @[Reg.scala 27:20]
  wire [1:0] _T_21245 = _T_22080 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21500 = _T_21499 | _T_21245; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_162; // @[Reg.scala 27:20]
  wire [1:0] _T_21246 = _T_22083 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21501 = _T_21500 | _T_21246; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_163; // @[Reg.scala 27:20]
  wire [1:0] _T_21247 = _T_22086 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21502 = _T_21501 | _T_21247; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_164; // @[Reg.scala 27:20]
  wire [1:0] _T_21248 = _T_22089 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21503 = _T_21502 | _T_21248; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_165; // @[Reg.scala 27:20]
  wire [1:0] _T_21249 = _T_22092 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21504 = _T_21503 | _T_21249; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_166; // @[Reg.scala 27:20]
  wire [1:0] _T_21250 = _T_22095 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21505 = _T_21504 | _T_21250; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_167; // @[Reg.scala 27:20]
  wire [1:0] _T_21251 = _T_22098 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21506 = _T_21505 | _T_21251; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_168; // @[Reg.scala 27:20]
  wire [1:0] _T_21252 = _T_22101 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21507 = _T_21506 | _T_21252; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_169; // @[Reg.scala 27:20]
  wire [1:0] _T_21253 = _T_22104 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21508 = _T_21507 | _T_21253; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_170; // @[Reg.scala 27:20]
  wire [1:0] _T_21254 = _T_22107 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21509 = _T_21508 | _T_21254; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_171; // @[Reg.scala 27:20]
  wire [1:0] _T_21255 = _T_22110 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21510 = _T_21509 | _T_21255; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_172; // @[Reg.scala 27:20]
  wire [1:0] _T_21256 = _T_22113 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21511 = _T_21510 | _T_21256; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_173; // @[Reg.scala 27:20]
  wire [1:0] _T_21257 = _T_22116 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21512 = _T_21511 | _T_21257; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_174; // @[Reg.scala 27:20]
  wire [1:0] _T_21258 = _T_22119 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21513 = _T_21512 | _T_21258; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_175; // @[Reg.scala 27:20]
  wire [1:0] _T_21259 = _T_22122 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21514 = _T_21513 | _T_21259; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_176; // @[Reg.scala 27:20]
  wire [1:0] _T_21260 = _T_22125 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21515 = _T_21514 | _T_21260; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_177; // @[Reg.scala 27:20]
  wire [1:0] _T_21261 = _T_22128 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21516 = _T_21515 | _T_21261; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_178; // @[Reg.scala 27:20]
  wire [1:0] _T_21262 = _T_22131 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21517 = _T_21516 | _T_21262; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_179; // @[Reg.scala 27:20]
  wire [1:0] _T_21263 = _T_22134 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21518 = _T_21517 | _T_21263; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_180; // @[Reg.scala 27:20]
  wire [1:0] _T_21264 = _T_22137 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21519 = _T_21518 | _T_21264; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_181; // @[Reg.scala 27:20]
  wire [1:0] _T_21265 = _T_22140 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21520 = _T_21519 | _T_21265; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_182; // @[Reg.scala 27:20]
  wire [1:0] _T_21266 = _T_22143 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21521 = _T_21520 | _T_21266; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_183; // @[Reg.scala 27:20]
  wire [1:0] _T_21267 = _T_22146 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21522 = _T_21521 | _T_21267; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_184; // @[Reg.scala 27:20]
  wire [1:0] _T_21268 = _T_22149 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21523 = _T_21522 | _T_21268; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_185; // @[Reg.scala 27:20]
  wire [1:0] _T_21269 = _T_22152 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21524 = _T_21523 | _T_21269; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_186; // @[Reg.scala 27:20]
  wire [1:0] _T_21270 = _T_22155 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21525 = _T_21524 | _T_21270; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_187; // @[Reg.scala 27:20]
  wire [1:0] _T_21271 = _T_22158 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21526 = _T_21525 | _T_21271; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_188; // @[Reg.scala 27:20]
  wire [1:0] _T_21272 = _T_22161 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21527 = _T_21526 | _T_21272; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_189; // @[Reg.scala 27:20]
  wire [1:0] _T_21273 = _T_22164 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21528 = _T_21527 | _T_21273; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_190; // @[Reg.scala 27:20]
  wire [1:0] _T_21274 = _T_22167 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21529 = _T_21528 | _T_21274; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_191; // @[Reg.scala 27:20]
  wire [1:0] _T_21275 = _T_22170 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21530 = _T_21529 | _T_21275; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_192; // @[Reg.scala 27:20]
  wire [1:0] _T_21276 = _T_22173 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21531 = _T_21530 | _T_21276; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_193; // @[Reg.scala 27:20]
  wire [1:0] _T_21277 = _T_22176 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21532 = _T_21531 | _T_21277; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_194; // @[Reg.scala 27:20]
  wire [1:0] _T_21278 = _T_22179 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21533 = _T_21532 | _T_21278; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_195; // @[Reg.scala 27:20]
  wire [1:0] _T_21279 = _T_22182 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21534 = _T_21533 | _T_21279; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_196; // @[Reg.scala 27:20]
  wire [1:0] _T_21280 = _T_22185 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21535 = _T_21534 | _T_21280; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_197; // @[Reg.scala 27:20]
  wire [1:0] _T_21281 = _T_22188 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21536 = _T_21535 | _T_21281; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_198; // @[Reg.scala 27:20]
  wire [1:0] _T_21282 = _T_22191 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21537 = _T_21536 | _T_21282; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_199; // @[Reg.scala 27:20]
  wire [1:0] _T_21283 = _T_22194 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21538 = _T_21537 | _T_21283; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_200; // @[Reg.scala 27:20]
  wire [1:0] _T_21284 = _T_22197 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21539 = _T_21538 | _T_21284; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_201; // @[Reg.scala 27:20]
  wire [1:0] _T_21285 = _T_22200 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21540 = _T_21539 | _T_21285; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_202; // @[Reg.scala 27:20]
  wire [1:0] _T_21286 = _T_22203 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21541 = _T_21540 | _T_21286; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_203; // @[Reg.scala 27:20]
  wire [1:0] _T_21287 = _T_22206 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21542 = _T_21541 | _T_21287; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_204; // @[Reg.scala 27:20]
  wire [1:0] _T_21288 = _T_22209 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21543 = _T_21542 | _T_21288; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_205; // @[Reg.scala 27:20]
  wire [1:0] _T_21289 = _T_22212 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21544 = _T_21543 | _T_21289; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_206; // @[Reg.scala 27:20]
  wire [1:0] _T_21290 = _T_22215 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21545 = _T_21544 | _T_21290; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_207; // @[Reg.scala 27:20]
  wire [1:0] _T_21291 = _T_22218 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21546 = _T_21545 | _T_21291; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_208; // @[Reg.scala 27:20]
  wire [1:0] _T_21292 = _T_22221 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21547 = _T_21546 | _T_21292; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_209; // @[Reg.scala 27:20]
  wire [1:0] _T_21293 = _T_22224 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21548 = _T_21547 | _T_21293; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_210; // @[Reg.scala 27:20]
  wire [1:0] _T_21294 = _T_22227 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21549 = _T_21548 | _T_21294; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_211; // @[Reg.scala 27:20]
  wire [1:0] _T_21295 = _T_22230 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21550 = _T_21549 | _T_21295; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_212; // @[Reg.scala 27:20]
  wire [1:0] _T_21296 = _T_22233 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21551 = _T_21550 | _T_21296; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_213; // @[Reg.scala 27:20]
  wire [1:0] _T_21297 = _T_22236 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21552 = _T_21551 | _T_21297; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_214; // @[Reg.scala 27:20]
  wire [1:0] _T_21298 = _T_22239 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21553 = _T_21552 | _T_21298; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_215; // @[Reg.scala 27:20]
  wire [1:0] _T_21299 = _T_22242 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21554 = _T_21553 | _T_21299; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_216; // @[Reg.scala 27:20]
  wire [1:0] _T_21300 = _T_22245 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21555 = _T_21554 | _T_21300; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_217; // @[Reg.scala 27:20]
  wire [1:0] _T_21301 = _T_22248 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21556 = _T_21555 | _T_21301; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_218; // @[Reg.scala 27:20]
  wire [1:0] _T_21302 = _T_22251 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21557 = _T_21556 | _T_21302; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_219; // @[Reg.scala 27:20]
  wire [1:0] _T_21303 = _T_22254 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21558 = _T_21557 | _T_21303; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_220; // @[Reg.scala 27:20]
  wire [1:0] _T_21304 = _T_22257 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21559 = _T_21558 | _T_21304; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_221; // @[Reg.scala 27:20]
  wire [1:0] _T_21305 = _T_22260 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21560 = _T_21559 | _T_21305; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_222; // @[Reg.scala 27:20]
  wire [1:0] _T_21306 = _T_22263 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21561 = _T_21560 | _T_21306; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_223; // @[Reg.scala 27:20]
  wire [1:0] _T_21307 = _T_22266 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21562 = _T_21561 | _T_21307; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_224; // @[Reg.scala 27:20]
  wire [1:0] _T_21308 = _T_22269 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21563 = _T_21562 | _T_21308; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_225; // @[Reg.scala 27:20]
  wire [1:0] _T_21309 = _T_22272 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21564 = _T_21563 | _T_21309; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_226; // @[Reg.scala 27:20]
  wire [1:0] _T_21310 = _T_22275 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21565 = _T_21564 | _T_21310; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_227; // @[Reg.scala 27:20]
  wire [1:0] _T_21311 = _T_22278 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21566 = _T_21565 | _T_21311; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_228; // @[Reg.scala 27:20]
  wire [1:0] _T_21312 = _T_22281 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21567 = _T_21566 | _T_21312; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_229; // @[Reg.scala 27:20]
  wire [1:0] _T_21313 = _T_22284 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21568 = _T_21567 | _T_21313; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_230; // @[Reg.scala 27:20]
  wire [1:0] _T_21314 = _T_22287 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21569 = _T_21568 | _T_21314; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_231; // @[Reg.scala 27:20]
  wire [1:0] _T_21315 = _T_22290 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21570 = _T_21569 | _T_21315; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_232; // @[Reg.scala 27:20]
  wire [1:0] _T_21316 = _T_22293 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21571 = _T_21570 | _T_21316; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_233; // @[Reg.scala 27:20]
  wire [1:0] _T_21317 = _T_22296 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21572 = _T_21571 | _T_21317; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_234; // @[Reg.scala 27:20]
  wire [1:0] _T_21318 = _T_22299 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21573 = _T_21572 | _T_21318; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_235; // @[Reg.scala 27:20]
  wire [1:0] _T_21319 = _T_22302 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21574 = _T_21573 | _T_21319; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_236; // @[Reg.scala 27:20]
  wire [1:0] _T_21320 = _T_22305 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21575 = _T_21574 | _T_21320; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_237; // @[Reg.scala 27:20]
  wire [1:0] _T_21321 = _T_22308 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21576 = _T_21575 | _T_21321; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_238; // @[Reg.scala 27:20]
  wire [1:0] _T_21322 = _T_22311 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21577 = _T_21576 | _T_21322; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_239; // @[Reg.scala 27:20]
  wire [1:0] _T_21323 = _T_22314 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21578 = _T_21577 | _T_21323; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_240; // @[Reg.scala 27:20]
  wire [1:0] _T_21324 = _T_22317 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21579 = _T_21578 | _T_21324; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_241; // @[Reg.scala 27:20]
  wire [1:0] _T_21325 = _T_22320 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21580 = _T_21579 | _T_21325; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_242; // @[Reg.scala 27:20]
  wire [1:0] _T_21326 = _T_22323 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21581 = _T_21580 | _T_21326; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_243; // @[Reg.scala 27:20]
  wire [1:0] _T_21327 = _T_22326 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21582 = _T_21581 | _T_21327; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_244; // @[Reg.scala 27:20]
  wire [1:0] _T_21328 = _T_22329 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21583 = _T_21582 | _T_21328; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_245; // @[Reg.scala 27:20]
  wire [1:0] _T_21329 = _T_22332 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21584 = _T_21583 | _T_21329; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_246; // @[Reg.scala 27:20]
  wire [1:0] _T_21330 = _T_22335 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21585 = _T_21584 | _T_21330; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_247; // @[Reg.scala 27:20]
  wire [1:0] _T_21331 = _T_22338 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21586 = _T_21585 | _T_21331; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_248; // @[Reg.scala 27:20]
  wire [1:0] _T_21332 = _T_22341 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21587 = _T_21586 | _T_21332; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_249; // @[Reg.scala 27:20]
  wire [1:0] _T_21333 = _T_22344 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21588 = _T_21587 | _T_21333; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_250; // @[Reg.scala 27:20]
  wire [1:0] _T_21334 = _T_22347 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21589 = _T_21588 | _T_21334; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_251; // @[Reg.scala 27:20]
  wire [1:0] _T_21335 = _T_22350 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21590 = _T_21589 | _T_21335; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_252; // @[Reg.scala 27:20]
  wire [1:0] _T_21336 = _T_22353 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21591 = _T_21590 | _T_21336; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_253; // @[Reg.scala 27:20]
  wire [1:0] _T_21337 = _T_22356 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21592 = _T_21591 | _T_21337; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_254; // @[Reg.scala 27:20]
  wire [1:0] _T_21338 = _T_22359 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21593 = _T_21592 | _T_21338; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_255; // @[Reg.scala 27:20]
  wire [1:0] _T_21339 = _T_22362 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_f = _T_21593 | _T_21339; // @[Mux.scala 27:72]
  wire [1:0] _T_250 = _T_143 ? bht_bank0_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_251 = io_ifc_fetch_addr_f[0] ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank0_rd_data_f = _T_250 | _T_251; // @[Mux.scala 27:72]
  wire  _T_268 = bht_force_taken_f[0] | bht_vbank0_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 251:45]
  wire  _T_270 = _T_268 & vwayhit_f[0]; // @[el2_ifu_bp_ctl.scala 251:72]
  wire [1:0] bht_dir_f = {_T_265,_T_270}; // @[Cat.scala 29:58]
  wire  _T_14 = ~bht_dir_f[0]; // @[el2_ifu_bp_ctl.scala 106:23]
  wire [1:0] btb_sel_f = {_T_14,bht_dir_f[0]}; // @[Cat.scala 29:58]
  wire [1:0] fetch_start_f = {io_ifc_fetch_addr_f[0],_T_143}; // @[Cat.scala 29:58]
  wire  _T_32 = io_exu_mp_btag == fetch_rd_tag_f; // @[el2_ifu_bp_ctl.scala 122:46]
  wire  _T_33 = _T_32 & exu_mp_valid; // @[el2_ifu_bp_ctl.scala 122:66]
  wire  _T_34 = _T_33 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 122:81]
  wire  _T_35 = io_exu_mp_index == btb_rd_addr_f; // @[el2_ifu_bp_ctl.scala 122:117]
  wire  fetch_mp_collision_f = _T_34 & _T_35; // @[el2_ifu_bp_ctl.scala 122:102]
  wire  _T_36 = io_exu_mp_btag == fetch_rd_tag_p1_f; // @[el2_ifu_bp_ctl.scala 123:49]
  wire  _T_37 = _T_36 & exu_mp_valid; // @[el2_ifu_bp_ctl.scala 123:72]
  wire  _T_38 = _T_37 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 123:87]
  wire  _T_39 = io_exu_mp_index == btb_rd_addr_p1_f; // @[el2_ifu_bp_ctl.scala 123:123]
  wire  fetch_mp_collision_p1_f = _T_38 & _T_39; // @[el2_ifu_bp_ctl.scala 123:108]
  reg  exu_mp_way_f; // @[el2_ifu_bp_ctl.scala 127:55]
  reg  exu_flush_final_d1; // @[el2_ifu_bp_ctl.scala 128:61]
  wire [255:0] mp_wrindex_dec = 256'h1 << io_exu_mp_index; // @[el2_ifu_bp_ctl.scala 181:28]
  wire [255:0] fetch_wrindex_dec = 256'h1 << btb_rd_addr_f; // @[el2_ifu_bp_ctl.scala 183:31]
  wire [255:0] fetch_wrindex_p1_dec = 256'h1 << btb_rd_addr_p1_f; // @[el2_ifu_bp_ctl.scala 185:34]
  wire [255:0] _T_149 = exu_mp_valid ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] mp_wrlru_b0 = mp_wrindex_dec & _T_149; // @[el2_ifu_bp_ctl.scala 187:36]
  wire  _T_165 = vwayhit_f[0] | vwayhit_f[1]; // @[el2_ifu_bp_ctl.scala 191:42]
  wire  _T_166 = _T_165 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 191:58]
  wire  lru_update_valid_f = _T_166 & _T; // @[el2_ifu_bp_ctl.scala 191:79]
  wire [255:0] _T_169 = lru_update_valid_f ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] fetch_wrlru_b0 = fetch_wrindex_dec & _T_169; // @[el2_ifu_bp_ctl.scala 193:42]
  wire [255:0] fetch_wrlru_p1_b0 = fetch_wrindex_p1_dec & _T_169; // @[el2_ifu_bp_ctl.scala 194:48]
  wire [255:0] _T_172 = ~mp_wrlru_b0; // @[el2_ifu_bp_ctl.scala 196:25]
  wire [255:0] _T_173 = ~fetch_wrlru_b0; // @[el2_ifu_bp_ctl.scala 196:40]
  wire [255:0] btb_lru_b0_hold = _T_172 & _T_173; // @[el2_ifu_bp_ctl.scala 196:38]
  wire  _T_175 = ~io_exu_mp_pkt_way; // @[el2_ifu_bp_ctl.scala 201:33]
  wire [255:0] _T_178 = _T_175 ? mp_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_179 = tag_match_way0_f ? fetch_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_180 = tag_match_way0_p1_f ? fetch_wrlru_p1_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_181 = _T_178 | _T_179; // @[Mux.scala 27:72]
  wire [255:0] _T_182 = _T_181 | _T_180; // @[Mux.scala 27:72]
  reg [255:0] btb_lru_b0_f; // @[Reg.scala 27:20]
  wire [255:0] _T_184 = btb_lru_b0_hold & btb_lru_b0_f; // @[el2_ifu_bp_ctl.scala 203:100]
  wire [255:0] btb_lru_b0_ns = _T_182 | _T_184; // @[el2_ifu_bp_ctl.scala 203:82]
  wire [255:0] _T_186 = fetch_wrindex_dec & btb_lru_b0_f; // @[el2_ifu_bp_ctl.scala 205:78]
  wire  _T_187 = |_T_186; // @[el2_ifu_bp_ctl.scala 205:94]
  wire  btb_lru_rd_f = fetch_mp_collision_f ? exu_mp_way_f : _T_187; // @[el2_ifu_bp_ctl.scala 205:25]
  wire [255:0] _T_189 = fetch_wrindex_p1_dec & btb_lru_b0_f; // @[el2_ifu_bp_ctl.scala 207:87]
  wire  _T_190 = |_T_189; // @[el2_ifu_bp_ctl.scala 207:103]
  wire  btb_lru_rd_p1_f = fetch_mp_collision_p1_f ? exu_mp_way_f : _T_190; // @[el2_ifu_bp_ctl.scala 207:28]
  wire [1:0] _T_193 = {btb_lru_rd_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_196 = {btb_lru_rd_p1_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_197 = _T_143 ? _T_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_198 = io_ifc_fetch_addr_f[0] ? _T_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] btb_vlru_rd_f = _T_197 | _T_198; // @[Mux.scala 27:72]
  wire [1:0] _T_207 = {tag_match_way1_expanded_p1_f[0],tag_match_way1_expanded_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_208 = _T_143 ? tag_match_way1_expanded_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_209 = io_ifc_fetch_addr_f[0] ? _T_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] tag_match_vway1_expanded_f = _T_208 | _T_209; // @[Mux.scala 27:72]
  wire [1:0] _T_211 = ~vwayhit_f; // @[el2_ifu_bp_ctl.scala 215:47]
  wire [1:0] _T_212 = _T_211 & btb_vlru_rd_f; // @[el2_ifu_bp_ctl.scala 215:58]
  wire  _T_213 = io_ifc_fetch_req_f | exu_mp_valid; // @[el2_ifu_bp_ctl.scala 217:75]
  wire [15:0] _T_228 = btb_sel_f[1] ? btb_vbank1_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_229 = btb_sel_f[0] ? btb_vbank0_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_230 = _T_228 | _T_229; // @[Mux.scala 27:72]
  wire [16:0] btb_sel_data_f = {{1'd0}, _T_230}; // @[el2_ifu_bp_ctl.scala 230:18]
  wire [11:0] btb_rd_tgt_f = btb_sel_data_f[15:4]; // @[el2_ifu_bp_ctl.scala 225:36]
  wire  btb_rd_pc4_f = btb_sel_data_f[3]; // @[el2_ifu_bp_ctl.scala 226:36]
  wire  btb_rd_call_f = btb_sel_data_f[1]; // @[el2_ifu_bp_ctl.scala 227:37]
  wire  btb_rd_ret_f = btb_sel_data_f[0]; // @[el2_ifu_bp_ctl.scala 228:36]
  wire [1:0] _T_278 = {bht_vbank1_rd_data_f[1],bht_vbank0_rd_data_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] hist1_raw = bht_force_taken_f | _T_278; // @[el2_ifu_bp_ctl.scala 256:34]
  wire [1:0] _T_232 = vwayhit_f & hist1_raw; // @[el2_ifu_bp_ctl.scala 233:39]
  wire  _T_233 = |_T_232; // @[el2_ifu_bp_ctl.scala 233:52]
  wire  _T_234 = _T_233 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 233:56]
  wire  _T_235 = ~leak_one_f_d1; // @[el2_ifu_bp_ctl.scala 233:79]
  wire  _T_236 = _T_234 & _T_235; // @[el2_ifu_bp_ctl.scala 233:77]
  wire  _T_237 = ~io_dec_tlu_bpred_disable; // @[el2_ifu_bp_ctl.scala 233:96]
  wire  _T_273 = io_ifu_bp_hit_taken_f & btb_sel_f[1]; // @[el2_ifu_bp_ctl.scala 253:51]
  wire  _T_274 = ~io_ifu_bp_hit_taken_f; // @[el2_ifu_bp_ctl.scala 253:69]
  wire  _T_284 = vwayhit_f[1] & btb_vbank1_rd_data_f[4]; // @[el2_ifu_bp_ctl.scala 260:34]
  wire  _T_287 = vwayhit_f[0] & btb_vbank0_rd_data_f[4]; // @[el2_ifu_bp_ctl.scala 261:34]
  wire  _T_290 = ~btb_vbank1_rd_data_f[2]; // @[el2_ifu_bp_ctl.scala 263:37]
  wire  _T_291 = vwayhit_f[1] & _T_290; // @[el2_ifu_bp_ctl.scala 263:35]
  wire  _T_293 = _T_291 & btb_vbank1_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 263:65]
  wire  _T_296 = ~btb_vbank0_rd_data_f[2]; // @[el2_ifu_bp_ctl.scala 264:37]
  wire  _T_297 = vwayhit_f[0] & _T_296; // @[el2_ifu_bp_ctl.scala 264:35]
  wire  _T_299 = _T_297 & btb_vbank0_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 264:65]
  wire [1:0] num_valids = vwayhit_f[1] + vwayhit_f[0]; // @[el2_ifu_bp_ctl.scala 267:35]
  wire [1:0] _T_302 = btb_sel_f & bht_dir_f; // @[el2_ifu_bp_ctl.scala 269:28]
  wire  final_h = |_T_302; // @[el2_ifu_bp_ctl.scala 269:41]
  wire  _T_303 = num_valids == 2'h2; // @[el2_ifu_bp_ctl.scala 273:41]
  wire [7:0] _T_307 = {fghr[5:0],1'h0,final_h}; // @[Cat.scala 29:58]
  wire  _T_308 = num_valids == 2'h1; // @[el2_ifu_bp_ctl.scala 274:41]
  wire [7:0] _T_311 = {fghr[6:0],final_h}; // @[Cat.scala 29:58]
  wire  _T_312 = num_valids == 2'h0; // @[el2_ifu_bp_ctl.scala 275:41]
  wire [7:0] _T_315 = _T_303 ? _T_307 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_316 = _T_308 ? _T_311 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_317 = _T_312 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_318 = _T_315 | _T_316; // @[Mux.scala 27:72]
  wire [7:0] merged_ghr = _T_318 | _T_317; // @[Mux.scala 27:72]
  wire  _T_321 = ~exu_flush_final_d1; // @[el2_ifu_bp_ctl.scala 280:27]
  wire  _T_322 = _T_321 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 280:47]
  wire  _T_323 = _T_322 & io_ic_hit_f; // @[el2_ifu_bp_ctl.scala 280:68]
  wire  _T_325 = _T_323 & _T_235; // @[el2_ifu_bp_ctl.scala 280:82]
  wire  _T_328 = io_ifc_fetch_req_f & io_ic_hit_f; // @[el2_ifu_bp_ctl.scala 281:70]
  wire  _T_330 = _T_328 & _T_235; // @[el2_ifu_bp_ctl.scala 281:84]
  wire  _T_331 = ~_T_330; // @[el2_ifu_bp_ctl.scala 281:49]
  wire  _T_332 = _T_321 & _T_331; // @[el2_ifu_bp_ctl.scala 281:47]
  wire [7:0] _T_334 = exu_flush_final_d1 ? io_exu_mp_fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_335 = _T_325 ? merged_ghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_336 = _T_332 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_337 = _T_334 | _T_335; // @[Mux.scala 27:72]
  wire [1:0] _T_341 = io_dec_tlu_bpred_disable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_342 = ~_T_341; // @[el2_ifu_bp_ctl.scala 292:36]
  wire  _T_346 = ~fetch_start_f[0]; // @[el2_ifu_bp_ctl.scala 295:36]
  wire  _T_347 = bht_dir_f[0] & _T_346; // @[el2_ifu_bp_ctl.scala 295:34]
  wire  _T_351 = _T_14 & fetch_start_f[0]; // @[el2_ifu_bp_ctl.scala 295:72]
  wire  _T_352 = _T_347 | _T_351; // @[el2_ifu_bp_ctl.scala 295:55]
  wire  _T_355 = bht_dir_f[0] & fetch_start_f[0]; // @[el2_ifu_bp_ctl.scala 296:19]
  wire  _T_360 = _T_14 & _T_346; // @[el2_ifu_bp_ctl.scala 296:56]
  wire  _T_361 = _T_355 | _T_360; // @[el2_ifu_bp_ctl.scala 296:39]
  wire [1:0] bloc_f = {_T_352,_T_361}; // @[Cat.scala 29:58]
  wire  _T_365 = _T_14 & io_ifc_fetch_addr_f[0]; // @[el2_ifu_bp_ctl.scala 298:35]
  wire  _T_366 = ~btb_rd_pc4_f; // @[el2_ifu_bp_ctl.scala 298:62]
  wire  use_fa_plus = _T_365 & _T_366; // @[el2_ifu_bp_ctl.scala 298:60]
  wire  _T_369 = fetch_start_f[0] & btb_sel_f[0]; // @[el2_ifu_bp_ctl.scala 300:44]
  wire  btb_fg_crossing_f = _T_369 & btb_rd_pc4_f; // @[el2_ifu_bp_ctl.scala 300:59]
  wire  bp_total_branch_offset_f = bloc_f[1] ^ btb_rd_pc4_f; // @[el2_ifu_bp_ctl.scala 301:43]
  wire  _T_372 = io_ifc_fetch_req_f & _T_274; // @[el2_ifu_bp_ctl.scala 303:87]
  wire  _T_373 = _T_372 & io_ic_hit_f; // @[el2_ifu_bp_ctl.scala 303:112]
  reg [30:0] ifc_fetch_adder_prior; // @[Reg.scala 27:20]
  wire  _T_377 = ~btb_fg_crossing_f; // @[el2_ifu_bp_ctl.scala 308:32]
  wire  _T_378 = ~use_fa_plus; // @[el2_ifu_bp_ctl.scala 308:53]
  wire  _T_379 = _T_377 & _T_378; // @[el2_ifu_bp_ctl.scala 308:51]
  wire [29:0] _T_382 = use_fa_plus ? fetch_addr_p1_f : 30'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_383 = btb_fg_crossing_f ? ifc_fetch_adder_prior : 31'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_384 = _T_379 ? io_ifc_fetch_addr_f[30:1] : 30'h0; // @[Mux.scala 27:72]
  wire [30:0] _GEN_1036 = {{1'd0}, _T_382}; // @[Mux.scala 27:72]
  wire [30:0] _T_385 = _GEN_1036 | _T_383; // @[Mux.scala 27:72]
  wire [30:0] _GEN_1037 = {{1'd0}, _T_384}; // @[Mux.scala 27:72]
  wire [30:0] adder_pc_in_f = _T_385 | _GEN_1037; // @[Mux.scala 27:72]
  wire [31:0] _T_389 = {adder_pc_in_f[29:0],bp_total_branch_offset_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_390 = {btb_rd_tgt_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_393 = _T_389[12:1] + _T_390[12:1]; // @[el2_lib.scala 201:31]
  wire [18:0] _T_396 = _T_389[31:13] + 19'h1; // @[el2_lib.scala 202:27]
  wire [18:0] _T_399 = _T_389[31:13] - 19'h1; // @[el2_lib.scala 203:27]
  wire  _T_402 = ~_T_393[12]; // @[el2_lib.scala 205:27]
  wire  _T_403 = _T_390[12] ^ _T_402; // @[el2_lib.scala 205:25]
  wire  _T_406 = ~_T_390[12]; // @[el2_lib.scala 206:8]
  wire  _T_408 = _T_406 & _T_393[12]; // @[el2_lib.scala 206:14]
  wire  _T_412 = _T_390[12] & _T_402; // @[el2_lib.scala 207:13]
  wire [18:0] _T_414 = _T_403 ? _T_389[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_415 = _T_408 ? _T_396 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_416 = _T_412 ? _T_399 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_417 = _T_414 | _T_415; // @[Mux.scala 27:72]
  wire [18:0] _T_418 = _T_417 | _T_416; // @[Mux.scala 27:72]
  wire [31:0] bp_btb_target_adder_f = {_T_418,_T_393[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_422 = ~btb_rd_call_f; // @[el2_ifu_bp_ctl.scala 315:49]
  wire  _T_423 = btb_rd_ret_f & _T_422; // @[el2_ifu_bp_ctl.scala 315:47]
  reg [31:0] rets_out_0; // @[Reg.scala 27:20]
  wire  _T_425 = _T_423 & rets_out_0[0]; // @[el2_ifu_bp_ctl.scala 315:64]
  wire [12:0] _T_436 = {11'h0,_T_366,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_439 = _T_389[12:1] + _T_436[12:1]; // @[el2_lib.scala 201:31]
  wire  _T_448 = ~_T_439[12]; // @[el2_lib.scala 205:27]
  wire  _T_449 = _T_436[12] ^ _T_448; // @[el2_lib.scala 205:25]
  wire  _T_452 = ~_T_436[12]; // @[el2_lib.scala 206:8]
  wire  _T_454 = _T_452 & _T_439[12]; // @[el2_lib.scala 206:14]
  wire  _T_458 = _T_436[12] & _T_448; // @[el2_lib.scala 207:13]
  wire [18:0] _T_460 = _T_449 ? _T_389[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_461 = _T_454 ? _T_396 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_462 = _T_458 ? _T_399 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_463 = _T_460 | _T_461; // @[Mux.scala 27:72]
  wire [18:0] _T_464 = _T_463 | _T_462; // @[Mux.scala 27:72]
  wire [31:0] bp_rs_call_target_f = {_T_464,_T_439[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_468 = ~btb_rd_ret_f; // @[el2_ifu_bp_ctl.scala 321:33]
  wire  _T_469 = btb_rd_call_f & _T_468; // @[el2_ifu_bp_ctl.scala 321:31]
  wire  rs_push = _T_469 & io_ifu_bp_hit_taken_f; // @[el2_ifu_bp_ctl.scala 321:47]
  wire  rs_pop = _T_423 & io_ifu_bp_hit_taken_f; // @[el2_ifu_bp_ctl.scala 322:46]
  wire  _T_472 = ~rs_push; // @[el2_ifu_bp_ctl.scala 323:17]
  wire  _T_473 = ~rs_pop; // @[el2_ifu_bp_ctl.scala 323:28]
  wire  rs_hold = _T_472 & _T_473; // @[el2_ifu_bp_ctl.scala 323:26]
  wire  rsenable_0 = ~rs_hold; // @[el2_ifu_bp_ctl.scala 325:60]
  wire  rsenable_1 = rs_push | rs_pop; // @[el2_ifu_bp_ctl.scala 325:119]
  wire [31:0] _T_476 = {bp_rs_call_target_f[31:1],1'h1}; // @[Cat.scala 29:58]
  wire [31:0] _T_478 = rs_push ? _T_476 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_1; // @[Reg.scala 27:20]
  wire [31:0] _T_479 = rs_pop ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_0 = _T_478 | _T_479; // @[Mux.scala 27:72]
  wire [31:0] _T_483 = rs_push ? rets_out_0 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_2; // @[Reg.scala 27:20]
  wire [31:0] _T_484 = rs_pop ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_1 = _T_483 | _T_484; // @[Mux.scala 27:72]
  wire [31:0] _T_488 = rs_push ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_3; // @[Reg.scala 27:20]
  wire [31:0] _T_489 = rs_pop ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_2 = _T_488 | _T_489; // @[Mux.scala 27:72]
  wire [31:0] _T_493 = rs_push ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_4; // @[Reg.scala 27:20]
  wire [31:0] _T_494 = rs_pop ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_3 = _T_493 | _T_494; // @[Mux.scala 27:72]
  wire [31:0] _T_498 = rs_push ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_5; // @[Reg.scala 27:20]
  wire [31:0] _T_499 = rs_pop ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_4 = _T_498 | _T_499; // @[Mux.scala 27:72]
  wire [31:0] _T_503 = rs_push ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_6; // @[Reg.scala 27:20]
  wire [31:0] _T_504 = rs_pop ? rets_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_5 = _T_503 | _T_504; // @[Mux.scala 27:72]
  wire [31:0] _T_508 = rs_push ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_7; // @[Reg.scala 27:20]
  wire [31:0] _T_509 = rs_pop ? rets_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_6 = _T_508 | _T_509; // @[Mux.scala 27:72]
  wire  _T_527 = ~dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 336:35]
  wire  btb_valid = exu_mp_valid & _T_527; // @[el2_ifu_bp_ctl.scala 336:32]
  wire  _T_528 = io_exu_mp_pkt_pcall | io_exu_mp_pkt_pja; // @[el2_ifu_bp_ctl.scala 339:89]
  wire  _T_529 = io_exu_mp_pkt_pret | io_exu_mp_pkt_pja; // @[el2_ifu_bp_ctl.scala 339:113]
  wire [21:0] btb_wr_data = {io_exu_mp_btag,io_exu_mp_pkt_toffset,io_exu_mp_pkt_pc4,io_exu_mp_pkt_boffset,_T_528,_T_529,btb_valid}; // @[Cat.scala 29:58]
  wire  exu_mp_valid_write = exu_mp_valid & io_exu_mp_pkt_ataken; // @[el2_ifu_bp_ctl.scala 340:41]
  wire  _T_536 = _T_175 & exu_mp_valid_write; // @[el2_ifu_bp_ctl.scala 342:39]
  wire  _T_538 = _T_536 & _T_527; // @[el2_ifu_bp_ctl.scala 342:60]
  wire  _T_539 = ~io_dec_tlu_br0_r_pkt_way; // @[el2_ifu_bp_ctl.scala 342:87]
  wire  _T_540 = _T_539 & dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 342:104]
  wire  btb_wr_en_way0 = _T_538 | _T_540; // @[el2_ifu_bp_ctl.scala 342:83]
  wire  _T_541 = io_exu_mp_pkt_way & exu_mp_valid_write; // @[el2_ifu_bp_ctl.scala 343:36]
  wire  _T_543 = _T_541 & _T_527; // @[el2_ifu_bp_ctl.scala 343:57]
  wire  _T_544 = io_dec_tlu_br0_r_pkt_way & dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 343:98]
  wire  btb_wr_en_way1 = _T_543 | _T_544; // @[el2_ifu_bp_ctl.scala 343:80]
  wire [7:0] btb_wr_addr = dec_tlu_error_wb ? {{1'd0}, btb_error_addr_wb} : io_exu_mp_index; // @[el2_ifu_bp_ctl.scala 345:24]
  wire  middle_of_bank = io_exu_mp_pkt_pc4 ^ io_exu_mp_pkt_boffset; // @[el2_ifu_bp_ctl.scala 346:35]
  wire  _T_546 = ~io_exu_mp_pkt_pcall; // @[el2_ifu_bp_ctl.scala 347:43]
  wire  _T_547 = exu_mp_valid & _T_546; // @[el2_ifu_bp_ctl.scala 347:41]
  wire  _T_548 = ~io_exu_mp_pkt_pret; // @[el2_ifu_bp_ctl.scala 347:58]
  wire  _T_549 = _T_547 & _T_548; // @[el2_ifu_bp_ctl.scala 347:56]
  wire  _T_550 = ~io_exu_mp_pkt_pja; // @[el2_ifu_bp_ctl.scala 347:72]
  wire  _T_551 = _T_549 & _T_550; // @[el2_ifu_bp_ctl.scala 347:70]
  wire [1:0] _T_553 = _T_551 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_554 = ~middle_of_bank; // @[el2_ifu_bp_ctl.scala 347:106]
  wire [1:0] _T_555 = {middle_of_bank,_T_554}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en0 = _T_553 & _T_555; // @[el2_ifu_bp_ctl.scala 347:84]
  wire [1:0] _T_557 = io_dec_tlu_br0_r_pkt_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_558 = ~io_dec_tlu_br0_r_pkt_middle; // @[el2_ifu_bp_ctl.scala 348:75]
  wire [1:0] _T_559 = {io_dec_tlu_br0_r_pkt_middle,_T_558}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en2 = _T_557 & _T_559; // @[el2_ifu_bp_ctl.scala 348:46]
  wire [9:0] _T_560 = {io_exu_mp_index,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] mp_hashed = _T_560[9:2] ^ io_exu_mp_eghr; // @[el2_lib.scala 191:35]
  wire [9:0] _T_563 = {io_exu_i0_br_index_r,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] br0_hashed_wb = _T_563[9:2] ^ io_exu_i0_br_fghr_r; // @[el2_lib.scala 191:35]
  wire  _T_572 = btb_wr_addr == 8'h0; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_573 = _T_572 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_575 = btb_wr_addr == 8'h1; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_576 = _T_575 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_578 = btb_wr_addr == 8'h2; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_579 = _T_578 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_581 = btb_wr_addr == 8'h3; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_582 = _T_581 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_584 = btb_wr_addr == 8'h4; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_585 = _T_584 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_587 = btb_wr_addr == 8'h5; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_588 = _T_587 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_590 = btb_wr_addr == 8'h6; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_591 = _T_590 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_593 = btb_wr_addr == 8'h7; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_594 = _T_593 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_596 = btb_wr_addr == 8'h8; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_597 = _T_596 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_599 = btb_wr_addr == 8'h9; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_600 = _T_599 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_602 = btb_wr_addr == 8'ha; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_603 = _T_602 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_605 = btb_wr_addr == 8'hb; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_606 = _T_605 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_608 = btb_wr_addr == 8'hc; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_609 = _T_608 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_611 = btb_wr_addr == 8'hd; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_612 = _T_611 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_614 = btb_wr_addr == 8'he; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_615 = _T_614 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_617 = btb_wr_addr == 8'hf; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_618 = _T_617 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_620 = btb_wr_addr == 8'h10; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_621 = _T_620 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_623 = btb_wr_addr == 8'h11; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_624 = _T_623 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_626 = btb_wr_addr == 8'h12; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_627 = _T_626 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_629 = btb_wr_addr == 8'h13; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_630 = _T_629 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_632 = btb_wr_addr == 8'h14; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_633 = _T_632 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_635 = btb_wr_addr == 8'h15; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_636 = _T_635 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_638 = btb_wr_addr == 8'h16; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_639 = _T_638 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_641 = btb_wr_addr == 8'h17; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_642 = _T_641 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_644 = btb_wr_addr == 8'h18; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_645 = _T_644 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_647 = btb_wr_addr == 8'h19; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_648 = _T_647 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_650 = btb_wr_addr == 8'h1a; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_651 = _T_650 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_653 = btb_wr_addr == 8'h1b; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_654 = _T_653 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_656 = btb_wr_addr == 8'h1c; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_657 = _T_656 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_659 = btb_wr_addr == 8'h1d; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_660 = _T_659 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_662 = btb_wr_addr == 8'h1e; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_663 = _T_662 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_665 = btb_wr_addr == 8'h1f; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_666 = _T_665 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_668 = btb_wr_addr == 8'h20; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_669 = _T_668 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_671 = btb_wr_addr == 8'h21; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_672 = _T_671 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_674 = btb_wr_addr == 8'h22; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_675 = _T_674 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_677 = btb_wr_addr == 8'h23; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_678 = _T_677 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_680 = btb_wr_addr == 8'h24; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_681 = _T_680 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_683 = btb_wr_addr == 8'h25; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_684 = _T_683 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_686 = btb_wr_addr == 8'h26; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_687 = _T_686 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_689 = btb_wr_addr == 8'h27; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_690 = _T_689 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_692 = btb_wr_addr == 8'h28; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_693 = _T_692 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_695 = btb_wr_addr == 8'h29; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_696 = _T_695 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_698 = btb_wr_addr == 8'h2a; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_699 = _T_698 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_701 = btb_wr_addr == 8'h2b; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_702 = _T_701 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_704 = btb_wr_addr == 8'h2c; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_705 = _T_704 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_707 = btb_wr_addr == 8'h2d; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_708 = _T_707 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_710 = btb_wr_addr == 8'h2e; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_711 = _T_710 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_713 = btb_wr_addr == 8'h2f; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_714 = _T_713 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_716 = btb_wr_addr == 8'h30; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_717 = _T_716 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_719 = btb_wr_addr == 8'h31; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_720 = _T_719 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_722 = btb_wr_addr == 8'h32; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_723 = _T_722 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_725 = btb_wr_addr == 8'h33; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_726 = _T_725 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_728 = btb_wr_addr == 8'h34; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_729 = _T_728 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_731 = btb_wr_addr == 8'h35; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_732 = _T_731 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_734 = btb_wr_addr == 8'h36; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_735 = _T_734 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_737 = btb_wr_addr == 8'h37; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_738 = _T_737 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_740 = btb_wr_addr == 8'h38; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_741 = _T_740 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_743 = btb_wr_addr == 8'h39; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_744 = _T_743 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_746 = btb_wr_addr == 8'h3a; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_747 = _T_746 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_749 = btb_wr_addr == 8'h3b; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_750 = _T_749 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_752 = btb_wr_addr == 8'h3c; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_753 = _T_752 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_755 = btb_wr_addr == 8'h3d; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_756 = _T_755 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_758 = btb_wr_addr == 8'h3e; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_759 = _T_758 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_761 = btb_wr_addr == 8'h3f; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_762 = _T_761 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_764 = btb_wr_addr == 8'h40; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_765 = _T_764 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_767 = btb_wr_addr == 8'h41; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_768 = _T_767 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_770 = btb_wr_addr == 8'h42; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_771 = _T_770 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_773 = btb_wr_addr == 8'h43; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_774 = _T_773 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_776 = btb_wr_addr == 8'h44; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_777 = _T_776 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_779 = btb_wr_addr == 8'h45; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_780 = _T_779 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_782 = btb_wr_addr == 8'h46; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_783 = _T_782 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_785 = btb_wr_addr == 8'h47; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_786 = _T_785 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_788 = btb_wr_addr == 8'h48; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_789 = _T_788 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_791 = btb_wr_addr == 8'h49; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_792 = _T_791 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_794 = btb_wr_addr == 8'h4a; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_795 = _T_794 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_797 = btb_wr_addr == 8'h4b; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_798 = _T_797 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_800 = btb_wr_addr == 8'h4c; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_801 = _T_800 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_803 = btb_wr_addr == 8'h4d; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_804 = _T_803 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_806 = btb_wr_addr == 8'h4e; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_807 = _T_806 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_809 = btb_wr_addr == 8'h4f; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_810 = _T_809 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_812 = btb_wr_addr == 8'h50; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_813 = _T_812 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_815 = btb_wr_addr == 8'h51; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_816 = _T_815 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_818 = btb_wr_addr == 8'h52; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_819 = _T_818 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_821 = btb_wr_addr == 8'h53; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_822 = _T_821 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_824 = btb_wr_addr == 8'h54; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_825 = _T_824 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_827 = btb_wr_addr == 8'h55; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_828 = _T_827 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_830 = btb_wr_addr == 8'h56; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_831 = _T_830 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_833 = btb_wr_addr == 8'h57; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_834 = _T_833 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_836 = btb_wr_addr == 8'h58; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_837 = _T_836 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_839 = btb_wr_addr == 8'h59; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_840 = _T_839 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_842 = btb_wr_addr == 8'h5a; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_843 = _T_842 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_845 = btb_wr_addr == 8'h5b; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_846 = _T_845 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_848 = btb_wr_addr == 8'h5c; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_849 = _T_848 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_851 = btb_wr_addr == 8'h5d; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_852 = _T_851 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_854 = btb_wr_addr == 8'h5e; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_855 = _T_854 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_857 = btb_wr_addr == 8'h5f; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_858 = _T_857 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_860 = btb_wr_addr == 8'h60; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_861 = _T_860 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_863 = btb_wr_addr == 8'h61; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_864 = _T_863 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_866 = btb_wr_addr == 8'h62; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_867 = _T_866 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_869 = btb_wr_addr == 8'h63; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_870 = _T_869 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_872 = btb_wr_addr == 8'h64; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_873 = _T_872 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_875 = btb_wr_addr == 8'h65; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_876 = _T_875 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_878 = btb_wr_addr == 8'h66; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_879 = _T_878 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_881 = btb_wr_addr == 8'h67; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_882 = _T_881 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_884 = btb_wr_addr == 8'h68; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_885 = _T_884 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_887 = btb_wr_addr == 8'h69; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_888 = _T_887 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_890 = btb_wr_addr == 8'h6a; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_891 = _T_890 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_893 = btb_wr_addr == 8'h6b; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_894 = _T_893 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_896 = btb_wr_addr == 8'h6c; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_897 = _T_896 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_899 = btb_wr_addr == 8'h6d; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_900 = _T_899 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_902 = btb_wr_addr == 8'h6e; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_903 = _T_902 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_905 = btb_wr_addr == 8'h6f; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_906 = _T_905 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_908 = btb_wr_addr == 8'h70; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_909 = _T_908 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_911 = btb_wr_addr == 8'h71; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_912 = _T_911 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_914 = btb_wr_addr == 8'h72; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_915 = _T_914 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_917 = btb_wr_addr == 8'h73; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_918 = _T_917 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_920 = btb_wr_addr == 8'h74; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_921 = _T_920 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_923 = btb_wr_addr == 8'h75; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_924 = _T_923 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_926 = btb_wr_addr == 8'h76; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_927 = _T_926 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_929 = btb_wr_addr == 8'h77; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_930 = _T_929 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_932 = btb_wr_addr == 8'h78; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_933 = _T_932 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_935 = btb_wr_addr == 8'h79; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_936 = _T_935 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_938 = btb_wr_addr == 8'h7a; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_939 = _T_938 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_941 = btb_wr_addr == 8'h7b; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_942 = _T_941 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_944 = btb_wr_addr == 8'h7c; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_945 = _T_944 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_947 = btb_wr_addr == 8'h7d; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_948 = _T_947 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_950 = btb_wr_addr == 8'h7e; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_951 = _T_950 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_953 = btb_wr_addr == 8'h7f; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_954 = _T_953 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_956 = btb_wr_addr == 8'h80; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_957 = _T_956 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_959 = btb_wr_addr == 8'h81; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_960 = _T_959 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_962 = btb_wr_addr == 8'h82; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_963 = _T_962 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_965 = btb_wr_addr == 8'h83; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_966 = _T_965 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_968 = btb_wr_addr == 8'h84; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_969 = _T_968 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_971 = btb_wr_addr == 8'h85; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_972 = _T_971 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_974 = btb_wr_addr == 8'h86; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_975 = _T_974 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_977 = btb_wr_addr == 8'h87; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_978 = _T_977 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_980 = btb_wr_addr == 8'h88; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_981 = _T_980 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_983 = btb_wr_addr == 8'h89; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_984 = _T_983 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_986 = btb_wr_addr == 8'h8a; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_987 = _T_986 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_989 = btb_wr_addr == 8'h8b; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_990 = _T_989 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_992 = btb_wr_addr == 8'h8c; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_993 = _T_992 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_995 = btb_wr_addr == 8'h8d; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_996 = _T_995 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_998 = btb_wr_addr == 8'h8e; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_999 = _T_998 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1001 = btb_wr_addr == 8'h8f; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1002 = _T_1001 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1004 = btb_wr_addr == 8'h90; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1005 = _T_1004 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1007 = btb_wr_addr == 8'h91; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1008 = _T_1007 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1010 = btb_wr_addr == 8'h92; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1011 = _T_1010 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1013 = btb_wr_addr == 8'h93; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1014 = _T_1013 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1016 = btb_wr_addr == 8'h94; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1017 = _T_1016 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1019 = btb_wr_addr == 8'h95; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1020 = _T_1019 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1022 = btb_wr_addr == 8'h96; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1023 = _T_1022 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1025 = btb_wr_addr == 8'h97; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1026 = _T_1025 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1028 = btb_wr_addr == 8'h98; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1029 = _T_1028 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1031 = btb_wr_addr == 8'h99; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1032 = _T_1031 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1034 = btb_wr_addr == 8'h9a; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1035 = _T_1034 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1037 = btb_wr_addr == 8'h9b; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1038 = _T_1037 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1040 = btb_wr_addr == 8'h9c; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1041 = _T_1040 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1043 = btb_wr_addr == 8'h9d; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1044 = _T_1043 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1046 = btb_wr_addr == 8'h9e; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1047 = _T_1046 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1049 = btb_wr_addr == 8'h9f; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1050 = _T_1049 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1052 = btb_wr_addr == 8'ha0; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1053 = _T_1052 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1055 = btb_wr_addr == 8'ha1; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1056 = _T_1055 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1058 = btb_wr_addr == 8'ha2; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1059 = _T_1058 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1061 = btb_wr_addr == 8'ha3; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1062 = _T_1061 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1064 = btb_wr_addr == 8'ha4; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1065 = _T_1064 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1067 = btb_wr_addr == 8'ha5; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1068 = _T_1067 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1070 = btb_wr_addr == 8'ha6; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1071 = _T_1070 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1073 = btb_wr_addr == 8'ha7; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1074 = _T_1073 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1076 = btb_wr_addr == 8'ha8; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1077 = _T_1076 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1079 = btb_wr_addr == 8'ha9; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1080 = _T_1079 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1082 = btb_wr_addr == 8'haa; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1083 = _T_1082 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1085 = btb_wr_addr == 8'hab; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1086 = _T_1085 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1088 = btb_wr_addr == 8'hac; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1089 = _T_1088 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1091 = btb_wr_addr == 8'had; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1092 = _T_1091 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1094 = btb_wr_addr == 8'hae; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1095 = _T_1094 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1097 = btb_wr_addr == 8'haf; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1098 = _T_1097 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1100 = btb_wr_addr == 8'hb0; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1101 = _T_1100 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1103 = btb_wr_addr == 8'hb1; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1104 = _T_1103 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1106 = btb_wr_addr == 8'hb2; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1107 = _T_1106 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1109 = btb_wr_addr == 8'hb3; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1110 = _T_1109 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1112 = btb_wr_addr == 8'hb4; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1113 = _T_1112 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1115 = btb_wr_addr == 8'hb5; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1116 = _T_1115 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1118 = btb_wr_addr == 8'hb6; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1119 = _T_1118 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1121 = btb_wr_addr == 8'hb7; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1122 = _T_1121 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1124 = btb_wr_addr == 8'hb8; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1125 = _T_1124 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1127 = btb_wr_addr == 8'hb9; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1128 = _T_1127 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1130 = btb_wr_addr == 8'hba; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1131 = _T_1130 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1133 = btb_wr_addr == 8'hbb; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1134 = _T_1133 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1136 = btb_wr_addr == 8'hbc; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1137 = _T_1136 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1139 = btb_wr_addr == 8'hbd; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1140 = _T_1139 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1142 = btb_wr_addr == 8'hbe; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1143 = _T_1142 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1145 = btb_wr_addr == 8'hbf; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1146 = _T_1145 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1148 = btb_wr_addr == 8'hc0; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1149 = _T_1148 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1151 = btb_wr_addr == 8'hc1; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1152 = _T_1151 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1154 = btb_wr_addr == 8'hc2; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1155 = _T_1154 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1157 = btb_wr_addr == 8'hc3; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1158 = _T_1157 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1160 = btb_wr_addr == 8'hc4; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1161 = _T_1160 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1163 = btb_wr_addr == 8'hc5; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1164 = _T_1163 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1166 = btb_wr_addr == 8'hc6; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1167 = _T_1166 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1169 = btb_wr_addr == 8'hc7; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1170 = _T_1169 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1172 = btb_wr_addr == 8'hc8; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1173 = _T_1172 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1175 = btb_wr_addr == 8'hc9; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1176 = _T_1175 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1178 = btb_wr_addr == 8'hca; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1179 = _T_1178 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1181 = btb_wr_addr == 8'hcb; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1182 = _T_1181 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1184 = btb_wr_addr == 8'hcc; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1185 = _T_1184 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1187 = btb_wr_addr == 8'hcd; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1188 = _T_1187 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1190 = btb_wr_addr == 8'hce; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1191 = _T_1190 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1193 = btb_wr_addr == 8'hcf; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1194 = _T_1193 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1196 = btb_wr_addr == 8'hd0; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1197 = _T_1196 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1199 = btb_wr_addr == 8'hd1; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1200 = _T_1199 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1202 = btb_wr_addr == 8'hd2; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1203 = _T_1202 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1205 = btb_wr_addr == 8'hd3; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1206 = _T_1205 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1208 = btb_wr_addr == 8'hd4; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1209 = _T_1208 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1211 = btb_wr_addr == 8'hd5; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1212 = _T_1211 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1214 = btb_wr_addr == 8'hd6; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1215 = _T_1214 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1217 = btb_wr_addr == 8'hd7; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1218 = _T_1217 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1220 = btb_wr_addr == 8'hd8; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1221 = _T_1220 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1223 = btb_wr_addr == 8'hd9; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1224 = _T_1223 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1226 = btb_wr_addr == 8'hda; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1227 = _T_1226 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1229 = btb_wr_addr == 8'hdb; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1230 = _T_1229 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1232 = btb_wr_addr == 8'hdc; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1233 = _T_1232 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1235 = btb_wr_addr == 8'hdd; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1236 = _T_1235 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1238 = btb_wr_addr == 8'hde; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1239 = _T_1238 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1241 = btb_wr_addr == 8'hdf; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1242 = _T_1241 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1244 = btb_wr_addr == 8'he0; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1245 = _T_1244 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1247 = btb_wr_addr == 8'he1; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1248 = _T_1247 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1250 = btb_wr_addr == 8'he2; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1251 = _T_1250 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1253 = btb_wr_addr == 8'he3; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1254 = _T_1253 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1256 = btb_wr_addr == 8'he4; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1257 = _T_1256 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1259 = btb_wr_addr == 8'he5; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1260 = _T_1259 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1262 = btb_wr_addr == 8'he6; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1263 = _T_1262 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1265 = btb_wr_addr == 8'he7; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1266 = _T_1265 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1268 = btb_wr_addr == 8'he8; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1269 = _T_1268 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1271 = btb_wr_addr == 8'he9; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1272 = _T_1271 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1274 = btb_wr_addr == 8'hea; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1275 = _T_1274 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1277 = btb_wr_addr == 8'heb; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1278 = _T_1277 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1280 = btb_wr_addr == 8'hec; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1281 = _T_1280 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1283 = btb_wr_addr == 8'hed; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1284 = _T_1283 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1286 = btb_wr_addr == 8'hee; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1287 = _T_1286 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1289 = btb_wr_addr == 8'hef; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1290 = _T_1289 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1292 = btb_wr_addr == 8'hf0; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1293 = _T_1292 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1295 = btb_wr_addr == 8'hf1; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1296 = _T_1295 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1298 = btb_wr_addr == 8'hf2; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1299 = _T_1298 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1301 = btb_wr_addr == 8'hf3; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1302 = _T_1301 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1304 = btb_wr_addr == 8'hf4; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1305 = _T_1304 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1307 = btb_wr_addr == 8'hf5; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1308 = _T_1307 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1310 = btb_wr_addr == 8'hf6; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1311 = _T_1310 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1313 = btb_wr_addr == 8'hf7; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1314 = _T_1313 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1316 = btb_wr_addr == 8'hf8; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1317 = _T_1316 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1319 = btb_wr_addr == 8'hf9; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1320 = _T_1319 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1322 = btb_wr_addr == 8'hfa; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1323 = _T_1322 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1325 = btb_wr_addr == 8'hfb; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1326 = _T_1325 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1328 = btb_wr_addr == 8'hfc; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1329 = _T_1328 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1331 = btb_wr_addr == 8'hfd; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1332 = _T_1331 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1334 = btb_wr_addr == 8'hfe; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1335 = _T_1334 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1337 = btb_wr_addr == 8'hff; // @[el2_ifu_bp_ctl.scala 365:101]
  wire  _T_1338 = _T_1337 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 365:109]
  wire  _T_1341 = _T_572 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1344 = _T_575 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1347 = _T_578 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1350 = _T_581 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1353 = _T_584 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1356 = _T_587 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1359 = _T_590 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1362 = _T_593 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1365 = _T_596 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1368 = _T_599 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1371 = _T_602 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1374 = _T_605 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1377 = _T_608 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1380 = _T_611 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1383 = _T_614 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1386 = _T_617 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1389 = _T_620 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1392 = _T_623 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1395 = _T_626 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1398 = _T_629 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1401 = _T_632 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1404 = _T_635 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1407 = _T_638 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1410 = _T_641 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1413 = _T_644 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1416 = _T_647 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1419 = _T_650 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1422 = _T_653 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1425 = _T_656 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1428 = _T_659 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1431 = _T_662 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1434 = _T_665 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1437 = _T_668 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1440 = _T_671 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1443 = _T_674 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1446 = _T_677 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1449 = _T_680 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1452 = _T_683 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1455 = _T_686 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1458 = _T_689 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1461 = _T_692 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1464 = _T_695 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1467 = _T_698 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1470 = _T_701 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1473 = _T_704 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1476 = _T_707 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1479 = _T_710 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1482 = _T_713 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1485 = _T_716 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1488 = _T_719 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1491 = _T_722 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1494 = _T_725 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1497 = _T_728 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1500 = _T_731 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1503 = _T_734 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1506 = _T_737 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1509 = _T_740 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1512 = _T_743 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1515 = _T_746 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1518 = _T_749 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1521 = _T_752 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1524 = _T_755 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1527 = _T_758 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1530 = _T_761 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1533 = _T_764 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1536 = _T_767 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1539 = _T_770 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1542 = _T_773 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1545 = _T_776 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1548 = _T_779 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1551 = _T_782 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1554 = _T_785 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1557 = _T_788 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1560 = _T_791 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1563 = _T_794 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1566 = _T_797 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1569 = _T_800 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1572 = _T_803 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1575 = _T_806 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1578 = _T_809 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1581 = _T_812 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1584 = _T_815 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1587 = _T_818 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1590 = _T_821 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1593 = _T_824 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1596 = _T_827 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1599 = _T_830 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1602 = _T_833 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1605 = _T_836 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1608 = _T_839 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1611 = _T_842 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1614 = _T_845 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1617 = _T_848 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1620 = _T_851 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1623 = _T_854 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1626 = _T_857 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1629 = _T_860 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1632 = _T_863 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1635 = _T_866 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1638 = _T_869 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1641 = _T_872 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1644 = _T_875 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1647 = _T_878 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1650 = _T_881 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1653 = _T_884 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1656 = _T_887 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1659 = _T_890 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1662 = _T_893 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1665 = _T_896 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1668 = _T_899 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1671 = _T_902 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1674 = _T_905 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1677 = _T_908 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1680 = _T_911 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1683 = _T_914 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1686 = _T_917 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1689 = _T_920 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1692 = _T_923 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1695 = _T_926 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1698 = _T_929 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1701 = _T_932 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1704 = _T_935 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1707 = _T_938 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1710 = _T_941 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1713 = _T_944 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1716 = _T_947 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1719 = _T_950 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1722 = _T_953 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1725 = _T_956 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1728 = _T_959 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1731 = _T_962 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1734 = _T_965 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1737 = _T_968 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1740 = _T_971 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1743 = _T_974 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1746 = _T_977 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1749 = _T_980 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1752 = _T_983 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1755 = _T_986 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1758 = _T_989 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1761 = _T_992 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1764 = _T_995 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1767 = _T_998 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1770 = _T_1001 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1773 = _T_1004 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1776 = _T_1007 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1779 = _T_1010 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1782 = _T_1013 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1785 = _T_1016 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1788 = _T_1019 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1791 = _T_1022 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1794 = _T_1025 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1797 = _T_1028 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1800 = _T_1031 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1803 = _T_1034 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1806 = _T_1037 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1809 = _T_1040 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1812 = _T_1043 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1815 = _T_1046 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1818 = _T_1049 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1821 = _T_1052 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1824 = _T_1055 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1827 = _T_1058 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1830 = _T_1061 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1833 = _T_1064 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1836 = _T_1067 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1839 = _T_1070 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1842 = _T_1073 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1845 = _T_1076 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1848 = _T_1079 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1851 = _T_1082 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1854 = _T_1085 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1857 = _T_1088 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1860 = _T_1091 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1863 = _T_1094 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1866 = _T_1097 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1869 = _T_1100 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1872 = _T_1103 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1875 = _T_1106 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1878 = _T_1109 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1881 = _T_1112 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1884 = _T_1115 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1887 = _T_1118 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1890 = _T_1121 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1893 = _T_1124 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1896 = _T_1127 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1899 = _T_1130 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1902 = _T_1133 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1905 = _T_1136 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1908 = _T_1139 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1911 = _T_1142 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1914 = _T_1145 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1917 = _T_1148 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1920 = _T_1151 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1923 = _T_1154 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1926 = _T_1157 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1929 = _T_1160 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1932 = _T_1163 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1935 = _T_1166 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1938 = _T_1169 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1941 = _T_1172 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1944 = _T_1175 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1947 = _T_1178 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1950 = _T_1181 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1953 = _T_1184 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1956 = _T_1187 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1959 = _T_1190 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1962 = _T_1193 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1965 = _T_1196 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1968 = _T_1199 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1971 = _T_1202 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1974 = _T_1205 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1977 = _T_1208 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1980 = _T_1211 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1983 = _T_1214 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1986 = _T_1217 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1989 = _T_1220 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1992 = _T_1223 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1995 = _T_1226 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1998 = _T_1229 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2001 = _T_1232 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2004 = _T_1235 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2007 = _T_1238 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2010 = _T_1241 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2013 = _T_1244 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2016 = _T_1247 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2019 = _T_1250 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2022 = _T_1253 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2025 = _T_1256 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2028 = _T_1259 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2031 = _T_1262 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2034 = _T_1265 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2037 = _T_1268 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2040 = _T_1271 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2043 = _T_1274 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2046 = _T_1277 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2049 = _T_1280 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2052 = _T_1283 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2055 = _T_1286 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2058 = _T_1289 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2061 = _T_1292 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2064 = _T_1295 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2067 = _T_1298 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2070 = _T_1301 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2073 = _T_1304 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2076 = _T_1307 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2079 = _T_1310 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2082 = _T_1313 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2085 = _T_1316 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2088 = _T_1319 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2091 = _T_1322 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2094 = _T_1325 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2097 = _T_1328 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2100 = _T_1331 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2103 = _T_1334 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_2106 = _T_1337 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_6494 = br0_hashed_wb[3:0] == 4'h0; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6495 = bht_wr_en2[0] & _T_6494; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6497 = ~br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_6498 = _T_6495 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6503 = br0_hashed_wb[3:0] == 4'h1; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6504 = bht_wr_en2[0] & _T_6503; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6507 = _T_6504 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6512 = br0_hashed_wb[3:0] == 4'h2; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6513 = bht_wr_en2[0] & _T_6512; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6516 = _T_6513 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6521 = br0_hashed_wb[3:0] == 4'h3; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6522 = bht_wr_en2[0] & _T_6521; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6525 = _T_6522 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6530 = br0_hashed_wb[3:0] == 4'h4; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6531 = bht_wr_en2[0] & _T_6530; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6534 = _T_6531 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6539 = br0_hashed_wb[3:0] == 4'h5; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6540 = bht_wr_en2[0] & _T_6539; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6543 = _T_6540 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6548 = br0_hashed_wb[3:0] == 4'h6; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6549 = bht_wr_en2[0] & _T_6548; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6552 = _T_6549 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6557 = br0_hashed_wb[3:0] == 4'h7; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6558 = bht_wr_en2[0] & _T_6557; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6561 = _T_6558 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6566 = br0_hashed_wb[3:0] == 4'h8; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6567 = bht_wr_en2[0] & _T_6566; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6570 = _T_6567 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6575 = br0_hashed_wb[3:0] == 4'h9; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6576 = bht_wr_en2[0] & _T_6575; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6579 = _T_6576 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6584 = br0_hashed_wb[3:0] == 4'ha; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6585 = bht_wr_en2[0] & _T_6584; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6588 = _T_6585 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6593 = br0_hashed_wb[3:0] == 4'hb; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6594 = bht_wr_en2[0] & _T_6593; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6597 = _T_6594 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6602 = br0_hashed_wb[3:0] == 4'hc; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6603 = bht_wr_en2[0] & _T_6602; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6606 = _T_6603 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6611 = br0_hashed_wb[3:0] == 4'hd; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6612 = bht_wr_en2[0] & _T_6611; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6615 = _T_6612 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6620 = br0_hashed_wb[3:0] == 4'he; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6621 = bht_wr_en2[0] & _T_6620; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6624 = _T_6621 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6629 = br0_hashed_wb[3:0] == 4'hf; // @[el2_ifu_bp_ctl.scala 381:74]
  wire  _T_6630 = bht_wr_en2[0] & _T_6629; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_6633 = _T_6630 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6642 = _T_6495 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6651 = _T_6504 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6660 = _T_6513 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6669 = _T_6522 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6678 = _T_6531 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6687 = _T_6540 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6696 = _T_6549 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6705 = _T_6558 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6714 = _T_6567 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6723 = _T_6576 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6732 = _T_6585 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6741 = _T_6594 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6750 = _T_6603 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6759 = _T_6612 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6768 = _T_6621 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6777 = _T_6630 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire [1:0] _GEN_1038 = {{1'd0}, br0_hashed_wb[4]}; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_6785 = _GEN_1038 == 2'h2; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_6786 = _T_6495 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6795 = _T_6504 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6804 = _T_6513 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6813 = _T_6522 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6822 = _T_6531 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6831 = _T_6540 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6840 = _T_6549 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6849 = _T_6558 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6858 = _T_6567 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6867 = _T_6576 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6876 = _T_6585 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6885 = _T_6594 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6894 = _T_6603 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6903 = _T_6612 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6912 = _T_6621 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6921 = _T_6630 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6929 = _GEN_1038 == 2'h3; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_6930 = _T_6495 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6939 = _T_6504 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6948 = _T_6513 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6957 = _T_6522 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6966 = _T_6531 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6975 = _T_6540 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6984 = _T_6549 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_6993 = _T_6558 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7002 = _T_6567 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7011 = _T_6576 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7020 = _T_6585 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7029 = _T_6594 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7038 = _T_6603 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7047 = _T_6612 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7056 = _T_6621 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7065 = _T_6630 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire [2:0] _GEN_1070 = {{2'd0}, br0_hashed_wb[4]}; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_7073 = _GEN_1070 == 3'h4; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_7074 = _T_6495 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7083 = _T_6504 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7092 = _T_6513 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7101 = _T_6522 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7110 = _T_6531 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7119 = _T_6540 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7128 = _T_6549 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7137 = _T_6558 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7146 = _T_6567 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7155 = _T_6576 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7164 = _T_6585 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7173 = _T_6594 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7182 = _T_6603 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7191 = _T_6612 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7200 = _T_6621 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7209 = _T_6630 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7217 = _GEN_1070 == 3'h5; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_7218 = _T_6495 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7227 = _T_6504 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7236 = _T_6513 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7245 = _T_6522 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7254 = _T_6531 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7263 = _T_6540 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7272 = _T_6549 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7281 = _T_6558 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7290 = _T_6567 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7299 = _T_6576 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7308 = _T_6585 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7317 = _T_6594 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7326 = _T_6603 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7335 = _T_6612 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7344 = _T_6621 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7353 = _T_6630 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7361 = _GEN_1070 == 3'h6; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_7362 = _T_6495 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7371 = _T_6504 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7380 = _T_6513 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7389 = _T_6522 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7398 = _T_6531 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7407 = _T_6540 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7416 = _T_6549 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7425 = _T_6558 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7434 = _T_6567 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7443 = _T_6576 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7452 = _T_6585 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7461 = _T_6594 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7470 = _T_6603 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7479 = _T_6612 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7488 = _T_6621 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7497 = _T_6630 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7505 = _GEN_1070 == 3'h7; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_7506 = _T_6495 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7515 = _T_6504 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7524 = _T_6513 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7533 = _T_6522 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7542 = _T_6531 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7551 = _T_6540 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7560 = _T_6549 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7569 = _T_6558 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7578 = _T_6567 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7587 = _T_6576 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7596 = _T_6585 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7605 = _T_6594 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7614 = _T_6603 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7623 = _T_6612 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7632 = _T_6621 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7641 = _T_6630 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire [3:0] _GEN_1134 = {{3'd0}, br0_hashed_wb[4]}; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_7649 = _GEN_1134 == 4'h8; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_7650 = _T_6495 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7659 = _T_6504 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7668 = _T_6513 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7677 = _T_6522 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7686 = _T_6531 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7695 = _T_6540 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7704 = _T_6549 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7713 = _T_6558 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7722 = _T_6567 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7731 = _T_6576 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7740 = _T_6585 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7749 = _T_6594 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7758 = _T_6603 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7767 = _T_6612 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7776 = _T_6621 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7785 = _T_6630 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7793 = _GEN_1134 == 4'h9; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_7794 = _T_6495 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7803 = _T_6504 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7812 = _T_6513 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7821 = _T_6522 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7830 = _T_6531 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7839 = _T_6540 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7848 = _T_6549 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7857 = _T_6558 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7866 = _T_6567 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7875 = _T_6576 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7884 = _T_6585 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7893 = _T_6594 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7902 = _T_6603 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7911 = _T_6612 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7920 = _T_6621 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7929 = _T_6630 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7937 = _GEN_1134 == 4'ha; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_7938 = _T_6495 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7947 = _T_6504 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7956 = _T_6513 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7965 = _T_6522 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7974 = _T_6531 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7983 = _T_6540 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_7992 = _T_6549 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8001 = _T_6558 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8010 = _T_6567 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8019 = _T_6576 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8028 = _T_6585 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8037 = _T_6594 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8046 = _T_6603 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8055 = _T_6612 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8064 = _T_6621 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8073 = _T_6630 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8081 = _GEN_1134 == 4'hb; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_8082 = _T_6495 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8091 = _T_6504 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8100 = _T_6513 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8109 = _T_6522 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8118 = _T_6531 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8127 = _T_6540 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8136 = _T_6549 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8145 = _T_6558 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8154 = _T_6567 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8163 = _T_6576 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8172 = _T_6585 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8181 = _T_6594 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8190 = _T_6603 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8199 = _T_6612 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8208 = _T_6621 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8217 = _T_6630 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8225 = _GEN_1134 == 4'hc; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_8226 = _T_6495 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8235 = _T_6504 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8244 = _T_6513 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8253 = _T_6522 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8262 = _T_6531 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8271 = _T_6540 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8280 = _T_6549 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8289 = _T_6558 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8298 = _T_6567 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8307 = _T_6576 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8316 = _T_6585 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8325 = _T_6594 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8334 = _T_6603 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8343 = _T_6612 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8352 = _T_6621 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8361 = _T_6630 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8369 = _GEN_1134 == 4'hd; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_8370 = _T_6495 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8379 = _T_6504 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8388 = _T_6513 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8397 = _T_6522 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8406 = _T_6531 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8415 = _T_6540 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8424 = _T_6549 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8433 = _T_6558 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8442 = _T_6567 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8451 = _T_6576 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8460 = _T_6585 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8469 = _T_6594 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8478 = _T_6603 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8487 = _T_6612 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8496 = _T_6621 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8505 = _T_6630 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8513 = _GEN_1134 == 4'he; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_8514 = _T_6495 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8523 = _T_6504 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8532 = _T_6513 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8541 = _T_6522 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8550 = _T_6531 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8559 = _T_6540 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8568 = _T_6549 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8577 = _T_6558 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8586 = _T_6567 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8595 = _T_6576 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8604 = _T_6585 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8613 = _T_6594 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8622 = _T_6603 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8631 = _T_6612 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8640 = _T_6621 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8649 = _T_6630 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8657 = _GEN_1134 == 4'hf; // @[el2_ifu_bp_ctl.scala 381:171]
  wire  _T_8658 = _T_6495 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8667 = _T_6504 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8676 = _T_6513 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8685 = _T_6522 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8694 = _T_6531 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8703 = _T_6540 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8712 = _T_6549 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8721 = _T_6558 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8730 = _T_6567 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8739 = _T_6576 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8748 = _T_6585 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8757 = _T_6594 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8766 = _T_6603 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8775 = _T_6612 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8784 = _T_6621 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8793 = _T_6630 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8799 = bht_wr_en2[1] & _T_6494; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8802 = _T_8799 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8808 = bht_wr_en2[1] & _T_6503; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8811 = _T_8808 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8817 = bht_wr_en2[1] & _T_6512; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8820 = _T_8817 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8826 = bht_wr_en2[1] & _T_6521; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8829 = _T_8826 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8835 = bht_wr_en2[1] & _T_6530; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8838 = _T_8835 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8844 = bht_wr_en2[1] & _T_6539; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8847 = _T_8844 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8853 = bht_wr_en2[1] & _T_6548; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8856 = _T_8853 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8862 = bht_wr_en2[1] & _T_6557; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8865 = _T_8862 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8871 = bht_wr_en2[1] & _T_6566; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8874 = _T_8871 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8880 = bht_wr_en2[1] & _T_6575; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8883 = _T_8880 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8889 = bht_wr_en2[1] & _T_6584; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8892 = _T_8889 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8898 = bht_wr_en2[1] & _T_6593; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8901 = _T_8898 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8907 = bht_wr_en2[1] & _T_6602; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8910 = _T_8907 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8916 = bht_wr_en2[1] & _T_6611; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8919 = _T_8916 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8925 = bht_wr_en2[1] & _T_6620; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8928 = _T_8925 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8934 = bht_wr_en2[1] & _T_6629; // @[el2_ifu_bp_ctl.scala 381:23]
  wire  _T_8937 = _T_8934 & _T_6497; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8946 = _T_8799 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8955 = _T_8808 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8964 = _T_8817 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8973 = _T_8826 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8982 = _T_8835 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_8991 = _T_8844 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9000 = _T_8853 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9009 = _T_8862 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9018 = _T_8871 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9027 = _T_8880 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9036 = _T_8889 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9045 = _T_8898 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9054 = _T_8907 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9063 = _T_8916 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9072 = _T_8925 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9081 = _T_8934 & br0_hashed_wb[4]; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9090 = _T_8799 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9099 = _T_8808 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9108 = _T_8817 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9117 = _T_8826 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9126 = _T_8835 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9135 = _T_8844 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9144 = _T_8853 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9153 = _T_8862 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9162 = _T_8871 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9171 = _T_8880 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9180 = _T_8889 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9189 = _T_8898 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9198 = _T_8907 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9207 = _T_8916 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9216 = _T_8925 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9225 = _T_8934 & _T_6785; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9234 = _T_8799 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9243 = _T_8808 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9252 = _T_8817 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9261 = _T_8826 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9270 = _T_8835 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9279 = _T_8844 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9288 = _T_8853 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9297 = _T_8862 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9306 = _T_8871 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9315 = _T_8880 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9324 = _T_8889 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9333 = _T_8898 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9342 = _T_8907 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9351 = _T_8916 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9360 = _T_8925 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9369 = _T_8934 & _T_6929; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9378 = _T_8799 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9387 = _T_8808 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9396 = _T_8817 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9405 = _T_8826 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9414 = _T_8835 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9423 = _T_8844 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9432 = _T_8853 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9441 = _T_8862 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9450 = _T_8871 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9459 = _T_8880 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9468 = _T_8889 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9477 = _T_8898 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9486 = _T_8907 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9495 = _T_8916 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9504 = _T_8925 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9513 = _T_8934 & _T_7073; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9522 = _T_8799 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9531 = _T_8808 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9540 = _T_8817 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9549 = _T_8826 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9558 = _T_8835 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9567 = _T_8844 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9576 = _T_8853 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9585 = _T_8862 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9594 = _T_8871 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9603 = _T_8880 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9612 = _T_8889 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9621 = _T_8898 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9630 = _T_8907 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9639 = _T_8916 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9648 = _T_8925 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9657 = _T_8934 & _T_7217; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9666 = _T_8799 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9675 = _T_8808 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9684 = _T_8817 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9693 = _T_8826 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9702 = _T_8835 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9711 = _T_8844 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9720 = _T_8853 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9729 = _T_8862 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9738 = _T_8871 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9747 = _T_8880 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9756 = _T_8889 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9765 = _T_8898 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9774 = _T_8907 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9783 = _T_8916 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9792 = _T_8925 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9801 = _T_8934 & _T_7361; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9810 = _T_8799 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9819 = _T_8808 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9828 = _T_8817 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9837 = _T_8826 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9846 = _T_8835 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9855 = _T_8844 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9864 = _T_8853 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9873 = _T_8862 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9882 = _T_8871 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9891 = _T_8880 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9900 = _T_8889 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9909 = _T_8898 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9918 = _T_8907 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9927 = _T_8916 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9936 = _T_8925 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9945 = _T_8934 & _T_7505; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9954 = _T_8799 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9963 = _T_8808 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9972 = _T_8817 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9981 = _T_8826 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9990 = _T_8835 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_9999 = _T_8844 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10008 = _T_8853 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10017 = _T_8862 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10026 = _T_8871 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10035 = _T_8880 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10044 = _T_8889 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10053 = _T_8898 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10062 = _T_8907 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10071 = _T_8916 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10080 = _T_8925 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10089 = _T_8934 & _T_7649; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10098 = _T_8799 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10107 = _T_8808 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10116 = _T_8817 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10125 = _T_8826 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10134 = _T_8835 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10143 = _T_8844 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10152 = _T_8853 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10161 = _T_8862 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10170 = _T_8871 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10179 = _T_8880 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10188 = _T_8889 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10197 = _T_8898 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10206 = _T_8907 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10215 = _T_8916 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10224 = _T_8925 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10233 = _T_8934 & _T_7793; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10242 = _T_8799 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10251 = _T_8808 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10260 = _T_8817 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10269 = _T_8826 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10278 = _T_8835 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10287 = _T_8844 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10296 = _T_8853 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10305 = _T_8862 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10314 = _T_8871 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10323 = _T_8880 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10332 = _T_8889 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10341 = _T_8898 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10350 = _T_8907 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10359 = _T_8916 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10368 = _T_8925 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10377 = _T_8934 & _T_7937; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10386 = _T_8799 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10395 = _T_8808 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10404 = _T_8817 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10413 = _T_8826 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10422 = _T_8835 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10431 = _T_8844 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10440 = _T_8853 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10449 = _T_8862 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10458 = _T_8871 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10467 = _T_8880 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10476 = _T_8889 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10485 = _T_8898 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10494 = _T_8907 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10503 = _T_8916 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10512 = _T_8925 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10521 = _T_8934 & _T_8081; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10530 = _T_8799 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10539 = _T_8808 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10548 = _T_8817 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10557 = _T_8826 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10566 = _T_8835 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10575 = _T_8844 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10584 = _T_8853 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10593 = _T_8862 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10602 = _T_8871 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10611 = _T_8880 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10620 = _T_8889 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10629 = _T_8898 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10638 = _T_8907 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10647 = _T_8916 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10656 = _T_8925 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10665 = _T_8934 & _T_8225; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10674 = _T_8799 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10683 = _T_8808 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10692 = _T_8817 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10701 = _T_8826 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10710 = _T_8835 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10719 = _T_8844 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10728 = _T_8853 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10737 = _T_8862 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10746 = _T_8871 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10755 = _T_8880 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10764 = _T_8889 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10773 = _T_8898 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10782 = _T_8907 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10791 = _T_8916 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10800 = _T_8925 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10809 = _T_8934 & _T_8369; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10818 = _T_8799 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10827 = _T_8808 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10836 = _T_8817 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10845 = _T_8826 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10854 = _T_8835 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10863 = _T_8844 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10872 = _T_8853 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10881 = _T_8862 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10890 = _T_8871 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10899 = _T_8880 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10908 = _T_8889 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10917 = _T_8898 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10926 = _T_8907 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10935 = _T_8916 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10944 = _T_8925 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10953 = _T_8934 & _T_8513; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10962 = _T_8799 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10971 = _T_8808 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10980 = _T_8817 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10989 = _T_8826 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_10998 = _T_8835 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11007 = _T_8844 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11016 = _T_8853 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11025 = _T_8862 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11034 = _T_8871 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11043 = _T_8880 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11052 = _T_8889 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11061 = _T_8898 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11070 = _T_8907 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11079 = _T_8916 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11088 = _T_8925 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11097 = _T_8934 & _T_8657; // @[el2_ifu_bp_ctl.scala 381:86]
  wire  _T_11102 = mp_hashed[3:0] == 4'h0; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11103 = bht_wr_en0[0] & _T_11102; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11105 = mp_hashed[7:4] == 4'h0; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_11107 = _T_11103 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11113 = br0_hashed_wb[7:4] == 4'h0; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_11115 = _T_6495 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_0 = _T_11107 | _T_11115; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11119 = mp_hashed[3:0] == 4'h1; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11120 = bht_wr_en0[0] & _T_11119; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11124 = _T_11120 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11132 = _T_6504 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_1 = _T_11124 | _T_11132; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11136 = mp_hashed[3:0] == 4'h2; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11137 = bht_wr_en0[0] & _T_11136; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11141 = _T_11137 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11149 = _T_6513 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_2 = _T_11141 | _T_11149; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11153 = mp_hashed[3:0] == 4'h3; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11154 = bht_wr_en0[0] & _T_11153; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11158 = _T_11154 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11166 = _T_6522 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_3 = _T_11158 | _T_11166; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11170 = mp_hashed[3:0] == 4'h4; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11171 = bht_wr_en0[0] & _T_11170; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11175 = _T_11171 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11183 = _T_6531 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_4 = _T_11175 | _T_11183; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11187 = mp_hashed[3:0] == 4'h5; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11188 = bht_wr_en0[0] & _T_11187; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11192 = _T_11188 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11200 = _T_6540 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_5 = _T_11192 | _T_11200; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11204 = mp_hashed[3:0] == 4'h6; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11205 = bht_wr_en0[0] & _T_11204; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11209 = _T_11205 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11217 = _T_6549 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_6 = _T_11209 | _T_11217; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11221 = mp_hashed[3:0] == 4'h7; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11222 = bht_wr_en0[0] & _T_11221; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11226 = _T_11222 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11234 = _T_6558 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_7 = _T_11226 | _T_11234; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11238 = mp_hashed[3:0] == 4'h8; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11239 = bht_wr_en0[0] & _T_11238; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11243 = _T_11239 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11251 = _T_6567 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_8 = _T_11243 | _T_11251; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11255 = mp_hashed[3:0] == 4'h9; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11256 = bht_wr_en0[0] & _T_11255; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11260 = _T_11256 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11268 = _T_6576 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_9 = _T_11260 | _T_11268; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11272 = mp_hashed[3:0] == 4'ha; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11273 = bht_wr_en0[0] & _T_11272; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11277 = _T_11273 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11285 = _T_6585 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_10 = _T_11277 | _T_11285; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11289 = mp_hashed[3:0] == 4'hb; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11290 = bht_wr_en0[0] & _T_11289; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11294 = _T_11290 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11302 = _T_6594 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_11 = _T_11294 | _T_11302; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11306 = mp_hashed[3:0] == 4'hc; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11307 = bht_wr_en0[0] & _T_11306; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11311 = _T_11307 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11319 = _T_6603 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_12 = _T_11311 | _T_11319; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11323 = mp_hashed[3:0] == 4'hd; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11324 = bht_wr_en0[0] & _T_11323; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11328 = _T_11324 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11336 = _T_6612 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_13 = _T_11328 | _T_11336; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11340 = mp_hashed[3:0] == 4'he; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11341 = bht_wr_en0[0] & _T_11340; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11345 = _T_11341 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11353 = _T_6621 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_14 = _T_11345 | _T_11353; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11357 = mp_hashed[3:0] == 4'hf; // @[el2_ifu_bp_ctl.scala 385:97]
  wire  _T_11358 = bht_wr_en0[0] & _T_11357; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_11362 = _T_11358 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11370 = _T_6630 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_0_15 = _T_11362 | _T_11370; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11377 = mp_hashed[7:4] == 4'h1; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_11379 = _T_11103 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11385 = br0_hashed_wb[7:4] == 4'h1; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_11387 = _T_6495 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_0 = _T_11379 | _T_11387; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11396 = _T_11120 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11404 = _T_6504 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_1 = _T_11396 | _T_11404; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11413 = _T_11137 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11421 = _T_6513 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_2 = _T_11413 | _T_11421; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11430 = _T_11154 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11438 = _T_6522 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_3 = _T_11430 | _T_11438; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11447 = _T_11171 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11455 = _T_6531 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_4 = _T_11447 | _T_11455; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11464 = _T_11188 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11472 = _T_6540 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_5 = _T_11464 | _T_11472; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11481 = _T_11205 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11489 = _T_6549 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_6 = _T_11481 | _T_11489; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11498 = _T_11222 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11506 = _T_6558 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_7 = _T_11498 | _T_11506; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11515 = _T_11239 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11523 = _T_6567 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_8 = _T_11515 | _T_11523; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11532 = _T_11256 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11540 = _T_6576 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_9 = _T_11532 | _T_11540; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11549 = _T_11273 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11557 = _T_6585 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_10 = _T_11549 | _T_11557; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11566 = _T_11290 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11574 = _T_6594 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_11 = _T_11566 | _T_11574; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11583 = _T_11307 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11591 = _T_6603 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_12 = _T_11583 | _T_11591; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11600 = _T_11324 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11608 = _T_6612 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_13 = _T_11600 | _T_11608; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11617 = _T_11341 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11625 = _T_6621 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_14 = _T_11617 | _T_11625; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11634 = _T_11358 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11642 = _T_6630 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_1_15 = _T_11634 | _T_11642; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11649 = mp_hashed[7:4] == 4'h2; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_11651 = _T_11103 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11657 = br0_hashed_wb[7:4] == 4'h2; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_11659 = _T_6495 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_0 = _T_11651 | _T_11659; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11668 = _T_11120 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11676 = _T_6504 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_1 = _T_11668 | _T_11676; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11685 = _T_11137 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11693 = _T_6513 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_2 = _T_11685 | _T_11693; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11702 = _T_11154 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11710 = _T_6522 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_3 = _T_11702 | _T_11710; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11719 = _T_11171 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11727 = _T_6531 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_4 = _T_11719 | _T_11727; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11736 = _T_11188 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11744 = _T_6540 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_5 = _T_11736 | _T_11744; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11753 = _T_11205 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11761 = _T_6549 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_6 = _T_11753 | _T_11761; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11770 = _T_11222 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11778 = _T_6558 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_7 = _T_11770 | _T_11778; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11787 = _T_11239 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11795 = _T_6567 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_8 = _T_11787 | _T_11795; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11804 = _T_11256 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11812 = _T_6576 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_9 = _T_11804 | _T_11812; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11821 = _T_11273 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11829 = _T_6585 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_10 = _T_11821 | _T_11829; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11838 = _T_11290 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11846 = _T_6594 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_11 = _T_11838 | _T_11846; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11855 = _T_11307 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11863 = _T_6603 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_12 = _T_11855 | _T_11863; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11872 = _T_11324 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11880 = _T_6612 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_13 = _T_11872 | _T_11880; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11889 = _T_11341 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11897 = _T_6621 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_14 = _T_11889 | _T_11897; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11906 = _T_11358 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11914 = _T_6630 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_2_15 = _T_11906 | _T_11914; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11921 = mp_hashed[7:4] == 4'h3; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_11923 = _T_11103 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11929 = br0_hashed_wb[7:4] == 4'h3; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_11931 = _T_6495 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_0 = _T_11923 | _T_11931; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11940 = _T_11120 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11948 = _T_6504 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_1 = _T_11940 | _T_11948; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11957 = _T_11137 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11965 = _T_6513 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_2 = _T_11957 | _T_11965; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11974 = _T_11154 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11982 = _T_6522 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_3 = _T_11974 | _T_11982; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_11991 = _T_11171 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_11999 = _T_6531 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_4 = _T_11991 | _T_11999; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12008 = _T_11188 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12016 = _T_6540 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_5 = _T_12008 | _T_12016; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12025 = _T_11205 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12033 = _T_6549 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_6 = _T_12025 | _T_12033; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12042 = _T_11222 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12050 = _T_6558 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_7 = _T_12042 | _T_12050; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12059 = _T_11239 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12067 = _T_6567 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_8 = _T_12059 | _T_12067; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12076 = _T_11256 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12084 = _T_6576 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_9 = _T_12076 | _T_12084; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12093 = _T_11273 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12101 = _T_6585 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_10 = _T_12093 | _T_12101; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12110 = _T_11290 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12118 = _T_6594 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_11 = _T_12110 | _T_12118; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12127 = _T_11307 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12135 = _T_6603 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_12 = _T_12127 | _T_12135; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12144 = _T_11324 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12152 = _T_6612 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_13 = _T_12144 | _T_12152; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12161 = _T_11341 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12169 = _T_6621 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_14 = _T_12161 | _T_12169; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12178 = _T_11358 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12186 = _T_6630 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_3_15 = _T_12178 | _T_12186; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12193 = mp_hashed[7:4] == 4'h4; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_12195 = _T_11103 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12201 = br0_hashed_wb[7:4] == 4'h4; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_12203 = _T_6495 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_0 = _T_12195 | _T_12203; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12212 = _T_11120 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12220 = _T_6504 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_1 = _T_12212 | _T_12220; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12229 = _T_11137 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12237 = _T_6513 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_2 = _T_12229 | _T_12237; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12246 = _T_11154 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12254 = _T_6522 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_3 = _T_12246 | _T_12254; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12263 = _T_11171 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12271 = _T_6531 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_4 = _T_12263 | _T_12271; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12280 = _T_11188 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12288 = _T_6540 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_5 = _T_12280 | _T_12288; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12297 = _T_11205 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12305 = _T_6549 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_6 = _T_12297 | _T_12305; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12314 = _T_11222 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12322 = _T_6558 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_7 = _T_12314 | _T_12322; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12331 = _T_11239 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12339 = _T_6567 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_8 = _T_12331 | _T_12339; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12348 = _T_11256 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12356 = _T_6576 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_9 = _T_12348 | _T_12356; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12365 = _T_11273 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12373 = _T_6585 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_10 = _T_12365 | _T_12373; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12382 = _T_11290 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12390 = _T_6594 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_11 = _T_12382 | _T_12390; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12399 = _T_11307 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12407 = _T_6603 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_12 = _T_12399 | _T_12407; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12416 = _T_11324 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12424 = _T_6612 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_13 = _T_12416 | _T_12424; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12433 = _T_11341 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12441 = _T_6621 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_14 = _T_12433 | _T_12441; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12450 = _T_11358 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12458 = _T_6630 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_4_15 = _T_12450 | _T_12458; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12465 = mp_hashed[7:4] == 4'h5; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_12467 = _T_11103 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12473 = br0_hashed_wb[7:4] == 4'h5; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_12475 = _T_6495 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_0 = _T_12467 | _T_12475; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12484 = _T_11120 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12492 = _T_6504 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_1 = _T_12484 | _T_12492; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12501 = _T_11137 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12509 = _T_6513 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_2 = _T_12501 | _T_12509; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12518 = _T_11154 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12526 = _T_6522 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_3 = _T_12518 | _T_12526; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12535 = _T_11171 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12543 = _T_6531 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_4 = _T_12535 | _T_12543; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12552 = _T_11188 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12560 = _T_6540 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_5 = _T_12552 | _T_12560; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12569 = _T_11205 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12577 = _T_6549 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_6 = _T_12569 | _T_12577; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12586 = _T_11222 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12594 = _T_6558 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_7 = _T_12586 | _T_12594; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12603 = _T_11239 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12611 = _T_6567 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_8 = _T_12603 | _T_12611; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12620 = _T_11256 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12628 = _T_6576 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_9 = _T_12620 | _T_12628; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12637 = _T_11273 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12645 = _T_6585 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_10 = _T_12637 | _T_12645; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12654 = _T_11290 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12662 = _T_6594 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_11 = _T_12654 | _T_12662; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12671 = _T_11307 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12679 = _T_6603 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_12 = _T_12671 | _T_12679; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12688 = _T_11324 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12696 = _T_6612 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_13 = _T_12688 | _T_12696; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12705 = _T_11341 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12713 = _T_6621 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_14 = _T_12705 | _T_12713; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12722 = _T_11358 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12730 = _T_6630 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_5_15 = _T_12722 | _T_12730; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12737 = mp_hashed[7:4] == 4'h6; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_12739 = _T_11103 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12745 = br0_hashed_wb[7:4] == 4'h6; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_12747 = _T_6495 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_0 = _T_12739 | _T_12747; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12756 = _T_11120 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12764 = _T_6504 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_1 = _T_12756 | _T_12764; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12773 = _T_11137 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12781 = _T_6513 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_2 = _T_12773 | _T_12781; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12790 = _T_11154 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12798 = _T_6522 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_3 = _T_12790 | _T_12798; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12807 = _T_11171 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12815 = _T_6531 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_4 = _T_12807 | _T_12815; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12824 = _T_11188 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12832 = _T_6540 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_5 = _T_12824 | _T_12832; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12841 = _T_11205 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12849 = _T_6549 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_6 = _T_12841 | _T_12849; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12858 = _T_11222 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12866 = _T_6558 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_7 = _T_12858 | _T_12866; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12875 = _T_11239 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12883 = _T_6567 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_8 = _T_12875 | _T_12883; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12892 = _T_11256 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12900 = _T_6576 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_9 = _T_12892 | _T_12900; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12909 = _T_11273 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12917 = _T_6585 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_10 = _T_12909 | _T_12917; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12926 = _T_11290 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12934 = _T_6594 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_11 = _T_12926 | _T_12934; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12943 = _T_11307 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12951 = _T_6603 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_12 = _T_12943 | _T_12951; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12960 = _T_11324 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12968 = _T_6612 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_13 = _T_12960 | _T_12968; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12977 = _T_11341 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_12985 = _T_6621 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_14 = _T_12977 | _T_12985; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_12994 = _T_11358 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13002 = _T_6630 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_6_15 = _T_12994 | _T_13002; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13009 = mp_hashed[7:4] == 4'h7; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_13011 = _T_11103 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13017 = br0_hashed_wb[7:4] == 4'h7; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_13019 = _T_6495 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_0 = _T_13011 | _T_13019; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13028 = _T_11120 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13036 = _T_6504 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_1 = _T_13028 | _T_13036; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13045 = _T_11137 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13053 = _T_6513 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_2 = _T_13045 | _T_13053; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13062 = _T_11154 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13070 = _T_6522 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_3 = _T_13062 | _T_13070; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13079 = _T_11171 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13087 = _T_6531 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_4 = _T_13079 | _T_13087; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13096 = _T_11188 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13104 = _T_6540 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_5 = _T_13096 | _T_13104; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13113 = _T_11205 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13121 = _T_6549 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_6 = _T_13113 | _T_13121; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13130 = _T_11222 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13138 = _T_6558 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_7 = _T_13130 | _T_13138; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13147 = _T_11239 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13155 = _T_6567 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_8 = _T_13147 | _T_13155; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13164 = _T_11256 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13172 = _T_6576 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_9 = _T_13164 | _T_13172; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13181 = _T_11273 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13189 = _T_6585 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_10 = _T_13181 | _T_13189; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13198 = _T_11290 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13206 = _T_6594 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_11 = _T_13198 | _T_13206; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13215 = _T_11307 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13223 = _T_6603 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_12 = _T_13215 | _T_13223; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13232 = _T_11324 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13240 = _T_6612 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_13 = _T_13232 | _T_13240; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13249 = _T_11341 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13257 = _T_6621 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_14 = _T_13249 | _T_13257; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13266 = _T_11358 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13274 = _T_6630 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_7_15 = _T_13266 | _T_13274; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13281 = mp_hashed[7:4] == 4'h8; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_13283 = _T_11103 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13289 = br0_hashed_wb[7:4] == 4'h8; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_13291 = _T_6495 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_0 = _T_13283 | _T_13291; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13300 = _T_11120 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13308 = _T_6504 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_1 = _T_13300 | _T_13308; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13317 = _T_11137 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13325 = _T_6513 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_2 = _T_13317 | _T_13325; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13334 = _T_11154 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13342 = _T_6522 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_3 = _T_13334 | _T_13342; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13351 = _T_11171 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13359 = _T_6531 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_4 = _T_13351 | _T_13359; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13368 = _T_11188 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13376 = _T_6540 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_5 = _T_13368 | _T_13376; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13385 = _T_11205 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13393 = _T_6549 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_6 = _T_13385 | _T_13393; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13402 = _T_11222 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13410 = _T_6558 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_7 = _T_13402 | _T_13410; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13419 = _T_11239 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13427 = _T_6567 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_8 = _T_13419 | _T_13427; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13436 = _T_11256 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13444 = _T_6576 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_9 = _T_13436 | _T_13444; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13453 = _T_11273 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13461 = _T_6585 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_10 = _T_13453 | _T_13461; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13470 = _T_11290 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13478 = _T_6594 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_11 = _T_13470 | _T_13478; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13487 = _T_11307 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13495 = _T_6603 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_12 = _T_13487 | _T_13495; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13504 = _T_11324 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13512 = _T_6612 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_13 = _T_13504 | _T_13512; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13521 = _T_11341 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13529 = _T_6621 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_14 = _T_13521 | _T_13529; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13538 = _T_11358 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13546 = _T_6630 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_8_15 = _T_13538 | _T_13546; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13553 = mp_hashed[7:4] == 4'h9; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_13555 = _T_11103 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13561 = br0_hashed_wb[7:4] == 4'h9; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_13563 = _T_6495 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_0 = _T_13555 | _T_13563; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13572 = _T_11120 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13580 = _T_6504 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_1 = _T_13572 | _T_13580; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13589 = _T_11137 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13597 = _T_6513 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_2 = _T_13589 | _T_13597; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13606 = _T_11154 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13614 = _T_6522 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_3 = _T_13606 | _T_13614; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13623 = _T_11171 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13631 = _T_6531 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_4 = _T_13623 | _T_13631; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13640 = _T_11188 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13648 = _T_6540 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_5 = _T_13640 | _T_13648; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13657 = _T_11205 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13665 = _T_6549 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_6 = _T_13657 | _T_13665; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13674 = _T_11222 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13682 = _T_6558 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_7 = _T_13674 | _T_13682; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13691 = _T_11239 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13699 = _T_6567 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_8 = _T_13691 | _T_13699; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13708 = _T_11256 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13716 = _T_6576 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_9 = _T_13708 | _T_13716; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13725 = _T_11273 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13733 = _T_6585 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_10 = _T_13725 | _T_13733; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13742 = _T_11290 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13750 = _T_6594 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_11 = _T_13742 | _T_13750; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13759 = _T_11307 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13767 = _T_6603 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_12 = _T_13759 | _T_13767; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13776 = _T_11324 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13784 = _T_6612 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_13 = _T_13776 | _T_13784; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13793 = _T_11341 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13801 = _T_6621 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_14 = _T_13793 | _T_13801; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13810 = _T_11358 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13818 = _T_6630 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_9_15 = _T_13810 | _T_13818; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13825 = mp_hashed[7:4] == 4'ha; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_13827 = _T_11103 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13833 = br0_hashed_wb[7:4] == 4'ha; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_13835 = _T_6495 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_0 = _T_13827 | _T_13835; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13844 = _T_11120 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13852 = _T_6504 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_1 = _T_13844 | _T_13852; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13861 = _T_11137 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13869 = _T_6513 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_2 = _T_13861 | _T_13869; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13878 = _T_11154 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13886 = _T_6522 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_3 = _T_13878 | _T_13886; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13895 = _T_11171 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13903 = _T_6531 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_4 = _T_13895 | _T_13903; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13912 = _T_11188 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13920 = _T_6540 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_5 = _T_13912 | _T_13920; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13929 = _T_11205 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13937 = _T_6549 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_6 = _T_13929 | _T_13937; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13946 = _T_11222 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13954 = _T_6558 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_7 = _T_13946 | _T_13954; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13963 = _T_11239 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13971 = _T_6567 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_8 = _T_13963 | _T_13971; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13980 = _T_11256 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_13988 = _T_6576 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_9 = _T_13980 | _T_13988; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_13997 = _T_11273 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14005 = _T_6585 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_10 = _T_13997 | _T_14005; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14014 = _T_11290 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14022 = _T_6594 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_11 = _T_14014 | _T_14022; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14031 = _T_11307 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14039 = _T_6603 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_12 = _T_14031 | _T_14039; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14048 = _T_11324 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14056 = _T_6612 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_13 = _T_14048 | _T_14056; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14065 = _T_11341 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14073 = _T_6621 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_14 = _T_14065 | _T_14073; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14082 = _T_11358 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14090 = _T_6630 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_10_15 = _T_14082 | _T_14090; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14097 = mp_hashed[7:4] == 4'hb; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_14099 = _T_11103 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14105 = br0_hashed_wb[7:4] == 4'hb; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_14107 = _T_6495 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_0 = _T_14099 | _T_14107; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14116 = _T_11120 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14124 = _T_6504 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_1 = _T_14116 | _T_14124; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14133 = _T_11137 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14141 = _T_6513 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_2 = _T_14133 | _T_14141; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14150 = _T_11154 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14158 = _T_6522 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_3 = _T_14150 | _T_14158; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14167 = _T_11171 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14175 = _T_6531 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_4 = _T_14167 | _T_14175; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14184 = _T_11188 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14192 = _T_6540 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_5 = _T_14184 | _T_14192; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14201 = _T_11205 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14209 = _T_6549 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_6 = _T_14201 | _T_14209; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14218 = _T_11222 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14226 = _T_6558 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_7 = _T_14218 | _T_14226; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14235 = _T_11239 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14243 = _T_6567 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_8 = _T_14235 | _T_14243; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14252 = _T_11256 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14260 = _T_6576 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_9 = _T_14252 | _T_14260; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14269 = _T_11273 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14277 = _T_6585 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_10 = _T_14269 | _T_14277; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14286 = _T_11290 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14294 = _T_6594 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_11 = _T_14286 | _T_14294; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14303 = _T_11307 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14311 = _T_6603 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_12 = _T_14303 | _T_14311; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14320 = _T_11324 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14328 = _T_6612 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_13 = _T_14320 | _T_14328; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14337 = _T_11341 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14345 = _T_6621 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_14 = _T_14337 | _T_14345; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14354 = _T_11358 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14362 = _T_6630 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_11_15 = _T_14354 | _T_14362; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14369 = mp_hashed[7:4] == 4'hc; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_14371 = _T_11103 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14377 = br0_hashed_wb[7:4] == 4'hc; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_14379 = _T_6495 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_0 = _T_14371 | _T_14379; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14388 = _T_11120 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14396 = _T_6504 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_1 = _T_14388 | _T_14396; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14405 = _T_11137 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14413 = _T_6513 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_2 = _T_14405 | _T_14413; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14422 = _T_11154 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14430 = _T_6522 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_3 = _T_14422 | _T_14430; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14439 = _T_11171 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14447 = _T_6531 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_4 = _T_14439 | _T_14447; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14456 = _T_11188 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14464 = _T_6540 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_5 = _T_14456 | _T_14464; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14473 = _T_11205 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14481 = _T_6549 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_6 = _T_14473 | _T_14481; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14490 = _T_11222 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14498 = _T_6558 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_7 = _T_14490 | _T_14498; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14507 = _T_11239 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14515 = _T_6567 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_8 = _T_14507 | _T_14515; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14524 = _T_11256 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14532 = _T_6576 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_9 = _T_14524 | _T_14532; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14541 = _T_11273 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14549 = _T_6585 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_10 = _T_14541 | _T_14549; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14558 = _T_11290 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14566 = _T_6594 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_11 = _T_14558 | _T_14566; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14575 = _T_11307 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14583 = _T_6603 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_12 = _T_14575 | _T_14583; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14592 = _T_11324 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14600 = _T_6612 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_13 = _T_14592 | _T_14600; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14609 = _T_11341 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14617 = _T_6621 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_14 = _T_14609 | _T_14617; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14626 = _T_11358 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14634 = _T_6630 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_12_15 = _T_14626 | _T_14634; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14641 = mp_hashed[7:4] == 4'hd; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_14643 = _T_11103 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14649 = br0_hashed_wb[7:4] == 4'hd; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_14651 = _T_6495 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_0 = _T_14643 | _T_14651; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14660 = _T_11120 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14668 = _T_6504 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_1 = _T_14660 | _T_14668; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14677 = _T_11137 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14685 = _T_6513 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_2 = _T_14677 | _T_14685; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14694 = _T_11154 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14702 = _T_6522 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_3 = _T_14694 | _T_14702; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14711 = _T_11171 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14719 = _T_6531 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_4 = _T_14711 | _T_14719; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14728 = _T_11188 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14736 = _T_6540 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_5 = _T_14728 | _T_14736; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14745 = _T_11205 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14753 = _T_6549 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_6 = _T_14745 | _T_14753; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14762 = _T_11222 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14770 = _T_6558 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_7 = _T_14762 | _T_14770; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14779 = _T_11239 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14787 = _T_6567 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_8 = _T_14779 | _T_14787; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14796 = _T_11256 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14804 = _T_6576 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_9 = _T_14796 | _T_14804; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14813 = _T_11273 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14821 = _T_6585 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_10 = _T_14813 | _T_14821; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14830 = _T_11290 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14838 = _T_6594 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_11 = _T_14830 | _T_14838; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14847 = _T_11307 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14855 = _T_6603 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_12 = _T_14847 | _T_14855; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14864 = _T_11324 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14872 = _T_6612 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_13 = _T_14864 | _T_14872; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14881 = _T_11341 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14889 = _T_6621 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_14 = _T_14881 | _T_14889; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14898 = _T_11358 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14906 = _T_6630 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_13_15 = _T_14898 | _T_14906; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14913 = mp_hashed[7:4] == 4'he; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_14915 = _T_11103 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14921 = br0_hashed_wb[7:4] == 4'he; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_14923 = _T_6495 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_0 = _T_14915 | _T_14923; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14932 = _T_11120 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14940 = _T_6504 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_1 = _T_14932 | _T_14940; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14949 = _T_11137 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14957 = _T_6513 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_2 = _T_14949 | _T_14957; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14966 = _T_11154 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14974 = _T_6522 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_3 = _T_14966 | _T_14974; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_14983 = _T_11171 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_14991 = _T_6531 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_4 = _T_14983 | _T_14991; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15000 = _T_11188 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15008 = _T_6540 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_5 = _T_15000 | _T_15008; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15017 = _T_11205 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15025 = _T_6549 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_6 = _T_15017 | _T_15025; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15034 = _T_11222 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15042 = _T_6558 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_7 = _T_15034 | _T_15042; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15051 = _T_11239 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15059 = _T_6567 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_8 = _T_15051 | _T_15059; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15068 = _T_11256 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15076 = _T_6576 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_9 = _T_15068 | _T_15076; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15085 = _T_11273 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15093 = _T_6585 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_10 = _T_15085 | _T_15093; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15102 = _T_11290 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15110 = _T_6594 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_11 = _T_15102 | _T_15110; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15119 = _T_11307 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15127 = _T_6603 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_12 = _T_15119 | _T_15127; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15136 = _T_11324 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15144 = _T_6612 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_13 = _T_15136 | _T_15144; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15153 = _T_11341 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15161 = _T_6621 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_14 = _T_15153 | _T_15161; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15170 = _T_11358 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15178 = _T_6630 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_14_15 = _T_15170 | _T_15178; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15185 = mp_hashed[7:4] == 4'hf; // @[el2_ifu_bp_ctl.scala 385:186]
  wire  _T_15187 = _T_11103 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15193 = br0_hashed_wb[7:4] == 4'hf; // @[el2_ifu_bp_ctl.scala 386:163]
  wire  _T_15195 = _T_6495 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_0 = _T_15187 | _T_15195; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15204 = _T_11120 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15212 = _T_6504 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_1 = _T_15204 | _T_15212; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15221 = _T_11137 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15229 = _T_6513 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_2 = _T_15221 | _T_15229; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15238 = _T_11154 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15246 = _T_6522 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_3 = _T_15238 | _T_15246; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15255 = _T_11171 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15263 = _T_6531 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_4 = _T_15255 | _T_15263; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15272 = _T_11188 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15280 = _T_6540 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_5 = _T_15272 | _T_15280; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15289 = _T_11205 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15297 = _T_6549 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_6 = _T_15289 | _T_15297; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15306 = _T_11222 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15314 = _T_6558 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_7 = _T_15306 | _T_15314; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15323 = _T_11239 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15331 = _T_6567 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_8 = _T_15323 | _T_15331; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15340 = _T_11256 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15348 = _T_6576 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_9 = _T_15340 | _T_15348; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15357 = _T_11273 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15365 = _T_6585 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_10 = _T_15357 | _T_15365; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15374 = _T_11290 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15382 = _T_6594 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_11 = _T_15374 | _T_15382; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15391 = _T_11307 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15399 = _T_6603 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_12 = _T_15391 | _T_15399; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15408 = _T_11324 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15416 = _T_6612 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_13 = _T_15408 | _T_15416; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15425 = _T_11341 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15433 = _T_6621 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_14 = _T_15425 | _T_15433; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15442 = _T_11358 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15450 = _T_6630 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_0_15_15 = _T_15442 | _T_15450; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15455 = bht_wr_en0[1] & _T_11102; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15459 = _T_15455 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15467 = _T_8799 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_0 = _T_15459 | _T_15467; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15472 = bht_wr_en0[1] & _T_11119; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15476 = _T_15472 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15484 = _T_8808 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_1 = _T_15476 | _T_15484; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15489 = bht_wr_en0[1] & _T_11136; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15493 = _T_15489 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15501 = _T_8817 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_2 = _T_15493 | _T_15501; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15506 = bht_wr_en0[1] & _T_11153; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15510 = _T_15506 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15518 = _T_8826 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_3 = _T_15510 | _T_15518; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15523 = bht_wr_en0[1] & _T_11170; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15527 = _T_15523 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15535 = _T_8835 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_4 = _T_15527 | _T_15535; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15540 = bht_wr_en0[1] & _T_11187; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15544 = _T_15540 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15552 = _T_8844 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_5 = _T_15544 | _T_15552; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15557 = bht_wr_en0[1] & _T_11204; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15561 = _T_15557 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15569 = _T_8853 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_6 = _T_15561 | _T_15569; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15574 = bht_wr_en0[1] & _T_11221; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15578 = _T_15574 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15586 = _T_8862 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_7 = _T_15578 | _T_15586; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15591 = bht_wr_en0[1] & _T_11238; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15595 = _T_15591 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15603 = _T_8871 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_8 = _T_15595 | _T_15603; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15608 = bht_wr_en0[1] & _T_11255; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15612 = _T_15608 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15620 = _T_8880 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_9 = _T_15612 | _T_15620; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15625 = bht_wr_en0[1] & _T_11272; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15629 = _T_15625 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15637 = _T_8889 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_10 = _T_15629 | _T_15637; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15642 = bht_wr_en0[1] & _T_11289; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15646 = _T_15642 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15654 = _T_8898 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_11 = _T_15646 | _T_15654; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15659 = bht_wr_en0[1] & _T_11306; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15663 = _T_15659 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15671 = _T_8907 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_12 = _T_15663 | _T_15671; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15676 = bht_wr_en0[1] & _T_11323; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15680 = _T_15676 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15688 = _T_8916 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_13 = _T_15680 | _T_15688; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15693 = bht_wr_en0[1] & _T_11340; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15697 = _T_15693 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15705 = _T_8925 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_14 = _T_15697 | _T_15705; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15710 = bht_wr_en0[1] & _T_11357; // @[el2_ifu_bp_ctl.scala 385:45]
  wire  _T_15714 = _T_15710 & _T_11105; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15722 = _T_8934 & _T_11113; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_0_15 = _T_15714 | _T_15722; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15731 = _T_15455 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15739 = _T_8799 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_0 = _T_15731 | _T_15739; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15748 = _T_15472 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15756 = _T_8808 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_1 = _T_15748 | _T_15756; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15765 = _T_15489 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15773 = _T_8817 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_2 = _T_15765 | _T_15773; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15782 = _T_15506 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15790 = _T_8826 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_3 = _T_15782 | _T_15790; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15799 = _T_15523 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15807 = _T_8835 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_4 = _T_15799 | _T_15807; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15816 = _T_15540 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15824 = _T_8844 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_5 = _T_15816 | _T_15824; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15833 = _T_15557 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15841 = _T_8853 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_6 = _T_15833 | _T_15841; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15850 = _T_15574 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15858 = _T_8862 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_7 = _T_15850 | _T_15858; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15867 = _T_15591 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15875 = _T_8871 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_8 = _T_15867 | _T_15875; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15884 = _T_15608 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15892 = _T_8880 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_9 = _T_15884 | _T_15892; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15901 = _T_15625 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15909 = _T_8889 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_10 = _T_15901 | _T_15909; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15918 = _T_15642 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15926 = _T_8898 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_11 = _T_15918 | _T_15926; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15935 = _T_15659 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15943 = _T_8907 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_12 = _T_15935 | _T_15943; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15952 = _T_15676 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15960 = _T_8916 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_13 = _T_15952 | _T_15960; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15969 = _T_15693 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15977 = _T_8925 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_14 = _T_15969 | _T_15977; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_15986 = _T_15710 & _T_11377; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_15994 = _T_8934 & _T_11385; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_1_15 = _T_15986 | _T_15994; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16003 = _T_15455 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16011 = _T_8799 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_0 = _T_16003 | _T_16011; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16020 = _T_15472 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16028 = _T_8808 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_1 = _T_16020 | _T_16028; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16037 = _T_15489 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16045 = _T_8817 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_2 = _T_16037 | _T_16045; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16054 = _T_15506 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16062 = _T_8826 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_3 = _T_16054 | _T_16062; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16071 = _T_15523 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16079 = _T_8835 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_4 = _T_16071 | _T_16079; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16088 = _T_15540 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16096 = _T_8844 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_5 = _T_16088 | _T_16096; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16105 = _T_15557 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16113 = _T_8853 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_6 = _T_16105 | _T_16113; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16122 = _T_15574 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16130 = _T_8862 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_7 = _T_16122 | _T_16130; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16139 = _T_15591 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16147 = _T_8871 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_8 = _T_16139 | _T_16147; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16156 = _T_15608 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16164 = _T_8880 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_9 = _T_16156 | _T_16164; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16173 = _T_15625 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16181 = _T_8889 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_10 = _T_16173 | _T_16181; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16190 = _T_15642 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16198 = _T_8898 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_11 = _T_16190 | _T_16198; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16207 = _T_15659 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16215 = _T_8907 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_12 = _T_16207 | _T_16215; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16224 = _T_15676 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16232 = _T_8916 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_13 = _T_16224 | _T_16232; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16241 = _T_15693 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16249 = _T_8925 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_14 = _T_16241 | _T_16249; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16258 = _T_15710 & _T_11649; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16266 = _T_8934 & _T_11657; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_2_15 = _T_16258 | _T_16266; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16275 = _T_15455 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16283 = _T_8799 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_0 = _T_16275 | _T_16283; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16292 = _T_15472 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16300 = _T_8808 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_1 = _T_16292 | _T_16300; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16309 = _T_15489 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16317 = _T_8817 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_2 = _T_16309 | _T_16317; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16326 = _T_15506 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16334 = _T_8826 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_3 = _T_16326 | _T_16334; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16343 = _T_15523 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16351 = _T_8835 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_4 = _T_16343 | _T_16351; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16360 = _T_15540 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16368 = _T_8844 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_5 = _T_16360 | _T_16368; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16377 = _T_15557 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16385 = _T_8853 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_6 = _T_16377 | _T_16385; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16394 = _T_15574 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16402 = _T_8862 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_7 = _T_16394 | _T_16402; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16411 = _T_15591 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16419 = _T_8871 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_8 = _T_16411 | _T_16419; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16428 = _T_15608 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16436 = _T_8880 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_9 = _T_16428 | _T_16436; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16445 = _T_15625 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16453 = _T_8889 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_10 = _T_16445 | _T_16453; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16462 = _T_15642 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16470 = _T_8898 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_11 = _T_16462 | _T_16470; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16479 = _T_15659 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16487 = _T_8907 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_12 = _T_16479 | _T_16487; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16496 = _T_15676 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16504 = _T_8916 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_13 = _T_16496 | _T_16504; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16513 = _T_15693 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16521 = _T_8925 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_14 = _T_16513 | _T_16521; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16530 = _T_15710 & _T_11921; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16538 = _T_8934 & _T_11929; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_3_15 = _T_16530 | _T_16538; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16547 = _T_15455 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16555 = _T_8799 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_0 = _T_16547 | _T_16555; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16564 = _T_15472 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16572 = _T_8808 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_1 = _T_16564 | _T_16572; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16581 = _T_15489 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16589 = _T_8817 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_2 = _T_16581 | _T_16589; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16598 = _T_15506 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16606 = _T_8826 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_3 = _T_16598 | _T_16606; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16615 = _T_15523 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16623 = _T_8835 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_4 = _T_16615 | _T_16623; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16632 = _T_15540 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16640 = _T_8844 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_5 = _T_16632 | _T_16640; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16649 = _T_15557 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16657 = _T_8853 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_6 = _T_16649 | _T_16657; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16666 = _T_15574 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16674 = _T_8862 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_7 = _T_16666 | _T_16674; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16683 = _T_15591 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16691 = _T_8871 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_8 = _T_16683 | _T_16691; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16700 = _T_15608 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16708 = _T_8880 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_9 = _T_16700 | _T_16708; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16717 = _T_15625 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16725 = _T_8889 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_10 = _T_16717 | _T_16725; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16734 = _T_15642 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16742 = _T_8898 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_11 = _T_16734 | _T_16742; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16751 = _T_15659 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16759 = _T_8907 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_12 = _T_16751 | _T_16759; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16768 = _T_15676 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16776 = _T_8916 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_13 = _T_16768 | _T_16776; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16785 = _T_15693 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16793 = _T_8925 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_14 = _T_16785 | _T_16793; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16802 = _T_15710 & _T_12193; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16810 = _T_8934 & _T_12201; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_4_15 = _T_16802 | _T_16810; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16819 = _T_15455 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16827 = _T_8799 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_0 = _T_16819 | _T_16827; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16836 = _T_15472 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16844 = _T_8808 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_1 = _T_16836 | _T_16844; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16853 = _T_15489 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16861 = _T_8817 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_2 = _T_16853 | _T_16861; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16870 = _T_15506 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16878 = _T_8826 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_3 = _T_16870 | _T_16878; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16887 = _T_15523 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16895 = _T_8835 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_4 = _T_16887 | _T_16895; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16904 = _T_15540 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16912 = _T_8844 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_5 = _T_16904 | _T_16912; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16921 = _T_15557 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16929 = _T_8853 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_6 = _T_16921 | _T_16929; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16938 = _T_15574 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16946 = _T_8862 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_7 = _T_16938 | _T_16946; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16955 = _T_15591 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16963 = _T_8871 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_8 = _T_16955 | _T_16963; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16972 = _T_15608 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16980 = _T_8880 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_9 = _T_16972 | _T_16980; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_16989 = _T_15625 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_16997 = _T_8889 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_10 = _T_16989 | _T_16997; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17006 = _T_15642 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17014 = _T_8898 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_11 = _T_17006 | _T_17014; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17023 = _T_15659 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17031 = _T_8907 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_12 = _T_17023 | _T_17031; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17040 = _T_15676 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17048 = _T_8916 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_13 = _T_17040 | _T_17048; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17057 = _T_15693 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17065 = _T_8925 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_14 = _T_17057 | _T_17065; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17074 = _T_15710 & _T_12465; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17082 = _T_8934 & _T_12473; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_5_15 = _T_17074 | _T_17082; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17091 = _T_15455 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17099 = _T_8799 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_0 = _T_17091 | _T_17099; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17108 = _T_15472 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17116 = _T_8808 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_1 = _T_17108 | _T_17116; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17125 = _T_15489 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17133 = _T_8817 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_2 = _T_17125 | _T_17133; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17142 = _T_15506 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17150 = _T_8826 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_3 = _T_17142 | _T_17150; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17159 = _T_15523 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17167 = _T_8835 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_4 = _T_17159 | _T_17167; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17176 = _T_15540 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17184 = _T_8844 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_5 = _T_17176 | _T_17184; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17193 = _T_15557 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17201 = _T_8853 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_6 = _T_17193 | _T_17201; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17210 = _T_15574 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17218 = _T_8862 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_7 = _T_17210 | _T_17218; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17227 = _T_15591 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17235 = _T_8871 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_8 = _T_17227 | _T_17235; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17244 = _T_15608 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17252 = _T_8880 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_9 = _T_17244 | _T_17252; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17261 = _T_15625 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17269 = _T_8889 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_10 = _T_17261 | _T_17269; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17278 = _T_15642 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17286 = _T_8898 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_11 = _T_17278 | _T_17286; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17295 = _T_15659 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17303 = _T_8907 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_12 = _T_17295 | _T_17303; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17312 = _T_15676 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17320 = _T_8916 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_13 = _T_17312 | _T_17320; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17329 = _T_15693 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17337 = _T_8925 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_14 = _T_17329 | _T_17337; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17346 = _T_15710 & _T_12737; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17354 = _T_8934 & _T_12745; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_6_15 = _T_17346 | _T_17354; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17363 = _T_15455 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17371 = _T_8799 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_0 = _T_17363 | _T_17371; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17380 = _T_15472 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17388 = _T_8808 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_1 = _T_17380 | _T_17388; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17397 = _T_15489 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17405 = _T_8817 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_2 = _T_17397 | _T_17405; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17414 = _T_15506 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17422 = _T_8826 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_3 = _T_17414 | _T_17422; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17431 = _T_15523 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17439 = _T_8835 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_4 = _T_17431 | _T_17439; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17448 = _T_15540 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17456 = _T_8844 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_5 = _T_17448 | _T_17456; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17465 = _T_15557 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17473 = _T_8853 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_6 = _T_17465 | _T_17473; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17482 = _T_15574 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17490 = _T_8862 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_7 = _T_17482 | _T_17490; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17499 = _T_15591 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17507 = _T_8871 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_8 = _T_17499 | _T_17507; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17516 = _T_15608 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17524 = _T_8880 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_9 = _T_17516 | _T_17524; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17533 = _T_15625 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17541 = _T_8889 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_10 = _T_17533 | _T_17541; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17550 = _T_15642 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17558 = _T_8898 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_11 = _T_17550 | _T_17558; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17567 = _T_15659 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17575 = _T_8907 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_12 = _T_17567 | _T_17575; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17584 = _T_15676 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17592 = _T_8916 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_13 = _T_17584 | _T_17592; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17601 = _T_15693 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17609 = _T_8925 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_14 = _T_17601 | _T_17609; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17618 = _T_15710 & _T_13009; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17626 = _T_8934 & _T_13017; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_7_15 = _T_17618 | _T_17626; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17635 = _T_15455 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17643 = _T_8799 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_0 = _T_17635 | _T_17643; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17652 = _T_15472 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17660 = _T_8808 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_1 = _T_17652 | _T_17660; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17669 = _T_15489 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17677 = _T_8817 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_2 = _T_17669 | _T_17677; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17686 = _T_15506 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17694 = _T_8826 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_3 = _T_17686 | _T_17694; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17703 = _T_15523 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17711 = _T_8835 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_4 = _T_17703 | _T_17711; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17720 = _T_15540 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17728 = _T_8844 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_5 = _T_17720 | _T_17728; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17737 = _T_15557 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17745 = _T_8853 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_6 = _T_17737 | _T_17745; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17754 = _T_15574 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17762 = _T_8862 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_7 = _T_17754 | _T_17762; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17771 = _T_15591 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17779 = _T_8871 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_8 = _T_17771 | _T_17779; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17788 = _T_15608 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17796 = _T_8880 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_9 = _T_17788 | _T_17796; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17805 = _T_15625 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17813 = _T_8889 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_10 = _T_17805 | _T_17813; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17822 = _T_15642 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17830 = _T_8898 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_11 = _T_17822 | _T_17830; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17839 = _T_15659 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17847 = _T_8907 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_12 = _T_17839 | _T_17847; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17856 = _T_15676 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17864 = _T_8916 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_13 = _T_17856 | _T_17864; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17873 = _T_15693 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17881 = _T_8925 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_14 = _T_17873 | _T_17881; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17890 = _T_15710 & _T_13281; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17898 = _T_8934 & _T_13289; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_8_15 = _T_17890 | _T_17898; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17907 = _T_15455 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17915 = _T_8799 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_0 = _T_17907 | _T_17915; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17924 = _T_15472 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17932 = _T_8808 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_1 = _T_17924 | _T_17932; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17941 = _T_15489 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17949 = _T_8817 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_2 = _T_17941 | _T_17949; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17958 = _T_15506 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17966 = _T_8826 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_3 = _T_17958 | _T_17966; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17975 = _T_15523 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_17983 = _T_8835 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_4 = _T_17975 | _T_17983; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_17992 = _T_15540 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18000 = _T_8844 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_5 = _T_17992 | _T_18000; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18009 = _T_15557 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18017 = _T_8853 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_6 = _T_18009 | _T_18017; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18026 = _T_15574 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18034 = _T_8862 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_7 = _T_18026 | _T_18034; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18043 = _T_15591 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18051 = _T_8871 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_8 = _T_18043 | _T_18051; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18060 = _T_15608 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18068 = _T_8880 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_9 = _T_18060 | _T_18068; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18077 = _T_15625 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18085 = _T_8889 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_10 = _T_18077 | _T_18085; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18094 = _T_15642 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18102 = _T_8898 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_11 = _T_18094 | _T_18102; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18111 = _T_15659 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18119 = _T_8907 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_12 = _T_18111 | _T_18119; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18128 = _T_15676 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18136 = _T_8916 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_13 = _T_18128 | _T_18136; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18145 = _T_15693 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18153 = _T_8925 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_14 = _T_18145 | _T_18153; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18162 = _T_15710 & _T_13553; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18170 = _T_8934 & _T_13561; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_9_15 = _T_18162 | _T_18170; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18179 = _T_15455 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18187 = _T_8799 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_0 = _T_18179 | _T_18187; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18196 = _T_15472 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18204 = _T_8808 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_1 = _T_18196 | _T_18204; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18213 = _T_15489 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18221 = _T_8817 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_2 = _T_18213 | _T_18221; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18230 = _T_15506 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18238 = _T_8826 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_3 = _T_18230 | _T_18238; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18247 = _T_15523 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18255 = _T_8835 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_4 = _T_18247 | _T_18255; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18264 = _T_15540 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18272 = _T_8844 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_5 = _T_18264 | _T_18272; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18281 = _T_15557 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18289 = _T_8853 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_6 = _T_18281 | _T_18289; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18298 = _T_15574 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18306 = _T_8862 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_7 = _T_18298 | _T_18306; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18315 = _T_15591 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18323 = _T_8871 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_8 = _T_18315 | _T_18323; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18332 = _T_15608 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18340 = _T_8880 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_9 = _T_18332 | _T_18340; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18349 = _T_15625 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18357 = _T_8889 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_10 = _T_18349 | _T_18357; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18366 = _T_15642 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18374 = _T_8898 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_11 = _T_18366 | _T_18374; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18383 = _T_15659 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18391 = _T_8907 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_12 = _T_18383 | _T_18391; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18400 = _T_15676 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18408 = _T_8916 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_13 = _T_18400 | _T_18408; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18417 = _T_15693 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18425 = _T_8925 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_14 = _T_18417 | _T_18425; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18434 = _T_15710 & _T_13825; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18442 = _T_8934 & _T_13833; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_10_15 = _T_18434 | _T_18442; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18451 = _T_15455 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18459 = _T_8799 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_0 = _T_18451 | _T_18459; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18468 = _T_15472 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18476 = _T_8808 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_1 = _T_18468 | _T_18476; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18485 = _T_15489 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18493 = _T_8817 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_2 = _T_18485 | _T_18493; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18502 = _T_15506 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18510 = _T_8826 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_3 = _T_18502 | _T_18510; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18519 = _T_15523 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18527 = _T_8835 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_4 = _T_18519 | _T_18527; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18536 = _T_15540 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18544 = _T_8844 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_5 = _T_18536 | _T_18544; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18553 = _T_15557 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18561 = _T_8853 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_6 = _T_18553 | _T_18561; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18570 = _T_15574 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18578 = _T_8862 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_7 = _T_18570 | _T_18578; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18587 = _T_15591 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18595 = _T_8871 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_8 = _T_18587 | _T_18595; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18604 = _T_15608 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18612 = _T_8880 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_9 = _T_18604 | _T_18612; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18621 = _T_15625 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18629 = _T_8889 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_10 = _T_18621 | _T_18629; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18638 = _T_15642 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18646 = _T_8898 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_11 = _T_18638 | _T_18646; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18655 = _T_15659 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18663 = _T_8907 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_12 = _T_18655 | _T_18663; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18672 = _T_15676 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18680 = _T_8916 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_13 = _T_18672 | _T_18680; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18689 = _T_15693 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18697 = _T_8925 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_14 = _T_18689 | _T_18697; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18706 = _T_15710 & _T_14097; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18714 = _T_8934 & _T_14105; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_11_15 = _T_18706 | _T_18714; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18723 = _T_15455 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18731 = _T_8799 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_0 = _T_18723 | _T_18731; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18740 = _T_15472 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18748 = _T_8808 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_1 = _T_18740 | _T_18748; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18757 = _T_15489 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18765 = _T_8817 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_2 = _T_18757 | _T_18765; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18774 = _T_15506 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18782 = _T_8826 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_3 = _T_18774 | _T_18782; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18791 = _T_15523 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18799 = _T_8835 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_4 = _T_18791 | _T_18799; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18808 = _T_15540 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18816 = _T_8844 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_5 = _T_18808 | _T_18816; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18825 = _T_15557 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18833 = _T_8853 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_6 = _T_18825 | _T_18833; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18842 = _T_15574 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18850 = _T_8862 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_7 = _T_18842 | _T_18850; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18859 = _T_15591 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18867 = _T_8871 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_8 = _T_18859 | _T_18867; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18876 = _T_15608 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18884 = _T_8880 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_9 = _T_18876 | _T_18884; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18893 = _T_15625 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18901 = _T_8889 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_10 = _T_18893 | _T_18901; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18910 = _T_15642 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18918 = _T_8898 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_11 = _T_18910 | _T_18918; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18927 = _T_15659 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18935 = _T_8907 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_12 = _T_18927 | _T_18935; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18944 = _T_15676 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18952 = _T_8916 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_13 = _T_18944 | _T_18952; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18961 = _T_15693 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18969 = _T_8925 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_14 = _T_18961 | _T_18969; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18978 = _T_15710 & _T_14369; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_18986 = _T_8934 & _T_14377; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_12_15 = _T_18978 | _T_18986; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_18995 = _T_15455 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19003 = _T_8799 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_0 = _T_18995 | _T_19003; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19012 = _T_15472 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19020 = _T_8808 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_1 = _T_19012 | _T_19020; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19029 = _T_15489 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19037 = _T_8817 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_2 = _T_19029 | _T_19037; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19046 = _T_15506 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19054 = _T_8826 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_3 = _T_19046 | _T_19054; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19063 = _T_15523 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19071 = _T_8835 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_4 = _T_19063 | _T_19071; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19080 = _T_15540 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19088 = _T_8844 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_5 = _T_19080 | _T_19088; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19097 = _T_15557 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19105 = _T_8853 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_6 = _T_19097 | _T_19105; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19114 = _T_15574 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19122 = _T_8862 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_7 = _T_19114 | _T_19122; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19131 = _T_15591 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19139 = _T_8871 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_8 = _T_19131 | _T_19139; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19148 = _T_15608 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19156 = _T_8880 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_9 = _T_19148 | _T_19156; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19165 = _T_15625 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19173 = _T_8889 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_10 = _T_19165 | _T_19173; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19182 = _T_15642 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19190 = _T_8898 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_11 = _T_19182 | _T_19190; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19199 = _T_15659 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19207 = _T_8907 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_12 = _T_19199 | _T_19207; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19216 = _T_15676 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19224 = _T_8916 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_13 = _T_19216 | _T_19224; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19233 = _T_15693 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19241 = _T_8925 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_14 = _T_19233 | _T_19241; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19250 = _T_15710 & _T_14641; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19258 = _T_8934 & _T_14649; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_13_15 = _T_19250 | _T_19258; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19267 = _T_15455 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19275 = _T_8799 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_0 = _T_19267 | _T_19275; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19284 = _T_15472 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19292 = _T_8808 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_1 = _T_19284 | _T_19292; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19301 = _T_15489 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19309 = _T_8817 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_2 = _T_19301 | _T_19309; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19318 = _T_15506 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19326 = _T_8826 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_3 = _T_19318 | _T_19326; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19335 = _T_15523 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19343 = _T_8835 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_4 = _T_19335 | _T_19343; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19352 = _T_15540 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19360 = _T_8844 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_5 = _T_19352 | _T_19360; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19369 = _T_15557 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19377 = _T_8853 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_6 = _T_19369 | _T_19377; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19386 = _T_15574 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19394 = _T_8862 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_7 = _T_19386 | _T_19394; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19403 = _T_15591 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19411 = _T_8871 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_8 = _T_19403 | _T_19411; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19420 = _T_15608 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19428 = _T_8880 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_9 = _T_19420 | _T_19428; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19437 = _T_15625 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19445 = _T_8889 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_10 = _T_19437 | _T_19445; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19454 = _T_15642 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19462 = _T_8898 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_11 = _T_19454 | _T_19462; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19471 = _T_15659 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19479 = _T_8907 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_12 = _T_19471 | _T_19479; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19488 = _T_15676 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19496 = _T_8916 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_13 = _T_19488 | _T_19496; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19505 = _T_15693 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19513 = _T_8925 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_14 = _T_19505 | _T_19513; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19522 = _T_15710 & _T_14913; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19530 = _T_8934 & _T_14921; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_14_15 = _T_19522 | _T_19530; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19539 = _T_15455 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19547 = _T_8799 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_0 = _T_19539 | _T_19547; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19556 = _T_15472 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19564 = _T_8808 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_1 = _T_19556 | _T_19564; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19573 = _T_15489 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19581 = _T_8817 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_2 = _T_19573 | _T_19581; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19590 = _T_15506 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19598 = _T_8826 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_3 = _T_19590 | _T_19598; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19607 = _T_15523 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19615 = _T_8835 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_4 = _T_19607 | _T_19615; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19624 = _T_15540 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19632 = _T_8844 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_5 = _T_19624 | _T_19632; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19641 = _T_15557 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19649 = _T_8853 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_6 = _T_19641 | _T_19649; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19658 = _T_15574 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19666 = _T_8862 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_7 = _T_19658 | _T_19666; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19675 = _T_15591 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19683 = _T_8871 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_8 = _T_19675 | _T_19683; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19692 = _T_15608 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19700 = _T_8880 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_9 = _T_19692 | _T_19700; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19709 = _T_15625 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19717 = _T_8889 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_10 = _T_19709 | _T_19717; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19726 = _T_15642 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19734 = _T_8898 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_11 = _T_19726 | _T_19734; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19743 = _T_15659 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19751 = _T_8907 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_12 = _T_19743 | _T_19751; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19760 = _T_15676 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19768 = _T_8916 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_13 = _T_19760 | _T_19768; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19777 = _T_15693 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19785 = _T_8925 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_14 = _T_19777 | _T_19785; // @[el2_ifu_bp_ctl.scala 385:223]
  wire  _T_19794 = _T_15710 & _T_15185; // @[el2_ifu_bp_ctl.scala 385:110]
  wire  _T_19802 = _T_8934 & _T_15193; // @[el2_ifu_bp_ctl.scala 386:87]
  wire  bht_bank_sel_1_15_15 = _T_19794 | _T_19802; // @[el2_ifu_bp_ctl.scala 385:223]
  assign io_ifu_bp_hit_taken_f = _T_236 & _T_237; // @[el2_ifu_bp_ctl.scala 233:25]
  assign io_ifu_bp_btb_target_f = _T_425 ? rets_out_0[31:1] : bp_btb_target_adder_f[31:1]; // @[el2_ifu_bp_ctl.scala 315:26]
  assign io_ifu_bp_inst_mask_f = _T_273 | _T_274; // @[el2_ifu_bp_ctl.scala 253:25]
  assign io_ifu_bp_fghr_f = fghr; // @[el2_ifu_bp_ctl.scala 285:20]
  assign io_ifu_bp_way_f = tag_match_vway1_expanded_f | _T_212; // @[el2_ifu_bp_ctl.scala 287:19]
  assign io_ifu_bp_ret_f = {_T_293,_T_299}; // @[el2_ifu_bp_ctl.scala 293:19]
  assign io_ifu_bp_hist1_f = bht_force_taken_f | _T_278; // @[el2_ifu_bp_ctl.scala 288:21]
  assign io_ifu_bp_hist0_f = {bht_vbank1_rd_data_f[0],bht_vbank0_rd_data_f[0]}; // @[el2_ifu_bp_ctl.scala 289:21]
  assign io_ifu_bp_pc4_f = {_T_284,_T_287}; // @[el2_ifu_bp_ctl.scala 290:19]
  assign io_ifu_bp_valid_f = vwayhit_f & _T_342; // @[el2_ifu_bp_ctl.scala 292:21]
  assign io_ifu_bp_poffset_f = btb_sel_data_f[15:4]; // @[el2_ifu_bp_ctl.scala 305:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  leak_one_f_d1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_0 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_1 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_2 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_3 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_4 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_5 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_6 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_7 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_8 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_9 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_10 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_11 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_12 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_13 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_14 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_15 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_16 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_17 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_18 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_19 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_20 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_21 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_22 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_23 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_24 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_25 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_26 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_27 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_28 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_29 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_30 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_31 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_32 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_33 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_34 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_35 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_36 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_37 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_38 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_39 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_40 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_41 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_42 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_43 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_44 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_45 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_46 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_47 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_48 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_49 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_50 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_51 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_52 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_53 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_54 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_55 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_56 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_57 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_58 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_59 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_60 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_61 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_62 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_63 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_64 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_65 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_66 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_67 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_68 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_69 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_70 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_71 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_72 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_73 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_74 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_75 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_76 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_77 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_78 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_79 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_80 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_81 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_82 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_83 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_84 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_85 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_86 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_87 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_88 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_89 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_90 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_91 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_92 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_93 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_94 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_95 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_96 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_97 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_98 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_99 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_100 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_101 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_102 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_103 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_104 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_105 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_106 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_107 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_108 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_109 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_110 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_111 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_112 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_113 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_114 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_115 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_116 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_117 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_118 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_119 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_120 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_121 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_122 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_123 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_124 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_125 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_126 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_127 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_128 = _RAND_129[21:0];
  _RAND_130 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_129 = _RAND_130[21:0];
  _RAND_131 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_130 = _RAND_131[21:0];
  _RAND_132 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_131 = _RAND_132[21:0];
  _RAND_133 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_132 = _RAND_133[21:0];
  _RAND_134 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_133 = _RAND_134[21:0];
  _RAND_135 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_134 = _RAND_135[21:0];
  _RAND_136 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_135 = _RAND_136[21:0];
  _RAND_137 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_136 = _RAND_137[21:0];
  _RAND_138 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_137 = _RAND_138[21:0];
  _RAND_139 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_138 = _RAND_139[21:0];
  _RAND_140 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_139 = _RAND_140[21:0];
  _RAND_141 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_140 = _RAND_141[21:0];
  _RAND_142 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_141 = _RAND_142[21:0];
  _RAND_143 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_142 = _RAND_143[21:0];
  _RAND_144 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_143 = _RAND_144[21:0];
  _RAND_145 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_144 = _RAND_145[21:0];
  _RAND_146 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_145 = _RAND_146[21:0];
  _RAND_147 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_146 = _RAND_147[21:0];
  _RAND_148 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_147 = _RAND_148[21:0];
  _RAND_149 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_148 = _RAND_149[21:0];
  _RAND_150 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_149 = _RAND_150[21:0];
  _RAND_151 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_150 = _RAND_151[21:0];
  _RAND_152 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_151 = _RAND_152[21:0];
  _RAND_153 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_152 = _RAND_153[21:0];
  _RAND_154 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_153 = _RAND_154[21:0];
  _RAND_155 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_154 = _RAND_155[21:0];
  _RAND_156 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_155 = _RAND_156[21:0];
  _RAND_157 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_156 = _RAND_157[21:0];
  _RAND_158 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_157 = _RAND_158[21:0];
  _RAND_159 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_158 = _RAND_159[21:0];
  _RAND_160 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_159 = _RAND_160[21:0];
  _RAND_161 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_160 = _RAND_161[21:0];
  _RAND_162 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_161 = _RAND_162[21:0];
  _RAND_163 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_162 = _RAND_163[21:0];
  _RAND_164 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_163 = _RAND_164[21:0];
  _RAND_165 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_164 = _RAND_165[21:0];
  _RAND_166 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_165 = _RAND_166[21:0];
  _RAND_167 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_166 = _RAND_167[21:0];
  _RAND_168 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_167 = _RAND_168[21:0];
  _RAND_169 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_168 = _RAND_169[21:0];
  _RAND_170 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_169 = _RAND_170[21:0];
  _RAND_171 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_170 = _RAND_171[21:0];
  _RAND_172 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_171 = _RAND_172[21:0];
  _RAND_173 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_172 = _RAND_173[21:0];
  _RAND_174 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_173 = _RAND_174[21:0];
  _RAND_175 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_174 = _RAND_175[21:0];
  _RAND_176 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_175 = _RAND_176[21:0];
  _RAND_177 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_176 = _RAND_177[21:0];
  _RAND_178 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_177 = _RAND_178[21:0];
  _RAND_179 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_178 = _RAND_179[21:0];
  _RAND_180 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_179 = _RAND_180[21:0];
  _RAND_181 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_180 = _RAND_181[21:0];
  _RAND_182 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_181 = _RAND_182[21:0];
  _RAND_183 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_182 = _RAND_183[21:0];
  _RAND_184 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_183 = _RAND_184[21:0];
  _RAND_185 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_184 = _RAND_185[21:0];
  _RAND_186 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_185 = _RAND_186[21:0];
  _RAND_187 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_186 = _RAND_187[21:0];
  _RAND_188 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_187 = _RAND_188[21:0];
  _RAND_189 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_188 = _RAND_189[21:0];
  _RAND_190 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_189 = _RAND_190[21:0];
  _RAND_191 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_190 = _RAND_191[21:0];
  _RAND_192 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_191 = _RAND_192[21:0];
  _RAND_193 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_192 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_193 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_194 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_195 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_196 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_197 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_198 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_199 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_200 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_201 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_202 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_203 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_204 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_205 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_206 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_207 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_208 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_209 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_210 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_211 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_212 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_213 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_214 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_215 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_216 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_217 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_218 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_219 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_220 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_221 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_222 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_223 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_224 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_225 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_226 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_227 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_228 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_229 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_230 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_231 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_232 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_233 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_234 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_235 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_236 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_237 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_238 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_239 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_240 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_241 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_242 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_243 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_244 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_245 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_246 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_247 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_248 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_249 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_250 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_251 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_252 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_253 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_254 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_255 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  dec_tlu_way_wb_f = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_0 = _RAND_258[21:0];
  _RAND_259 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_1 = _RAND_259[21:0];
  _RAND_260 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_2 = _RAND_260[21:0];
  _RAND_261 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_3 = _RAND_261[21:0];
  _RAND_262 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_4 = _RAND_262[21:0];
  _RAND_263 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_5 = _RAND_263[21:0];
  _RAND_264 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_6 = _RAND_264[21:0];
  _RAND_265 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_7 = _RAND_265[21:0];
  _RAND_266 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_8 = _RAND_266[21:0];
  _RAND_267 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_9 = _RAND_267[21:0];
  _RAND_268 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_10 = _RAND_268[21:0];
  _RAND_269 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_11 = _RAND_269[21:0];
  _RAND_270 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_12 = _RAND_270[21:0];
  _RAND_271 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_13 = _RAND_271[21:0];
  _RAND_272 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_14 = _RAND_272[21:0];
  _RAND_273 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_15 = _RAND_273[21:0];
  _RAND_274 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_16 = _RAND_274[21:0];
  _RAND_275 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_17 = _RAND_275[21:0];
  _RAND_276 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_18 = _RAND_276[21:0];
  _RAND_277 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_19 = _RAND_277[21:0];
  _RAND_278 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_20 = _RAND_278[21:0];
  _RAND_279 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_21 = _RAND_279[21:0];
  _RAND_280 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_22 = _RAND_280[21:0];
  _RAND_281 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_23 = _RAND_281[21:0];
  _RAND_282 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_24 = _RAND_282[21:0];
  _RAND_283 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_25 = _RAND_283[21:0];
  _RAND_284 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_26 = _RAND_284[21:0];
  _RAND_285 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_27 = _RAND_285[21:0];
  _RAND_286 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_28 = _RAND_286[21:0];
  _RAND_287 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_29 = _RAND_287[21:0];
  _RAND_288 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_30 = _RAND_288[21:0];
  _RAND_289 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_31 = _RAND_289[21:0];
  _RAND_290 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_32 = _RAND_290[21:0];
  _RAND_291 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_33 = _RAND_291[21:0];
  _RAND_292 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_34 = _RAND_292[21:0];
  _RAND_293 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_35 = _RAND_293[21:0];
  _RAND_294 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_36 = _RAND_294[21:0];
  _RAND_295 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_37 = _RAND_295[21:0];
  _RAND_296 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_38 = _RAND_296[21:0];
  _RAND_297 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_39 = _RAND_297[21:0];
  _RAND_298 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_40 = _RAND_298[21:0];
  _RAND_299 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_41 = _RAND_299[21:0];
  _RAND_300 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_42 = _RAND_300[21:0];
  _RAND_301 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_43 = _RAND_301[21:0];
  _RAND_302 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_44 = _RAND_302[21:0];
  _RAND_303 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_45 = _RAND_303[21:0];
  _RAND_304 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_46 = _RAND_304[21:0];
  _RAND_305 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_47 = _RAND_305[21:0];
  _RAND_306 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_48 = _RAND_306[21:0];
  _RAND_307 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_49 = _RAND_307[21:0];
  _RAND_308 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_50 = _RAND_308[21:0];
  _RAND_309 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_51 = _RAND_309[21:0];
  _RAND_310 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_52 = _RAND_310[21:0];
  _RAND_311 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_53 = _RAND_311[21:0];
  _RAND_312 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_54 = _RAND_312[21:0];
  _RAND_313 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_55 = _RAND_313[21:0];
  _RAND_314 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_56 = _RAND_314[21:0];
  _RAND_315 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_57 = _RAND_315[21:0];
  _RAND_316 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_58 = _RAND_316[21:0];
  _RAND_317 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_59 = _RAND_317[21:0];
  _RAND_318 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_60 = _RAND_318[21:0];
  _RAND_319 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_61 = _RAND_319[21:0];
  _RAND_320 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_62 = _RAND_320[21:0];
  _RAND_321 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_63 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_64 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_65 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_66 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_67 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_68 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_69 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_70 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_71 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_72 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_73 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_74 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_75 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_76 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_77 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_78 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_79 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_80 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_81 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_82 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_83 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_84 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_85 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_86 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_87 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_88 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_89 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_90 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_91 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_92 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_93 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_94 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_95 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_96 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_97 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_98 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_99 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_100 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_101 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_102 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_103 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_104 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_105 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_106 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_107 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_108 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_109 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_110 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_111 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_112 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_113 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_114 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_115 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_116 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_117 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_118 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_119 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_120 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_121 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_122 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_123 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_124 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_125 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_126 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_127 = _RAND_385[21:0];
  _RAND_386 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_128 = _RAND_386[21:0];
  _RAND_387 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_129 = _RAND_387[21:0];
  _RAND_388 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_130 = _RAND_388[21:0];
  _RAND_389 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_131 = _RAND_389[21:0];
  _RAND_390 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_132 = _RAND_390[21:0];
  _RAND_391 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_133 = _RAND_391[21:0];
  _RAND_392 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_134 = _RAND_392[21:0];
  _RAND_393 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_135 = _RAND_393[21:0];
  _RAND_394 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_136 = _RAND_394[21:0];
  _RAND_395 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_137 = _RAND_395[21:0];
  _RAND_396 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_138 = _RAND_396[21:0];
  _RAND_397 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_139 = _RAND_397[21:0];
  _RAND_398 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_140 = _RAND_398[21:0];
  _RAND_399 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_141 = _RAND_399[21:0];
  _RAND_400 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_142 = _RAND_400[21:0];
  _RAND_401 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_143 = _RAND_401[21:0];
  _RAND_402 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_144 = _RAND_402[21:0];
  _RAND_403 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_145 = _RAND_403[21:0];
  _RAND_404 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_146 = _RAND_404[21:0];
  _RAND_405 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_147 = _RAND_405[21:0];
  _RAND_406 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_148 = _RAND_406[21:0];
  _RAND_407 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_149 = _RAND_407[21:0];
  _RAND_408 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_150 = _RAND_408[21:0];
  _RAND_409 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_151 = _RAND_409[21:0];
  _RAND_410 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_152 = _RAND_410[21:0];
  _RAND_411 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_153 = _RAND_411[21:0];
  _RAND_412 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_154 = _RAND_412[21:0];
  _RAND_413 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_155 = _RAND_413[21:0];
  _RAND_414 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_156 = _RAND_414[21:0];
  _RAND_415 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_157 = _RAND_415[21:0];
  _RAND_416 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_158 = _RAND_416[21:0];
  _RAND_417 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_159 = _RAND_417[21:0];
  _RAND_418 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_160 = _RAND_418[21:0];
  _RAND_419 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_161 = _RAND_419[21:0];
  _RAND_420 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_162 = _RAND_420[21:0];
  _RAND_421 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_163 = _RAND_421[21:0];
  _RAND_422 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_164 = _RAND_422[21:0];
  _RAND_423 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_165 = _RAND_423[21:0];
  _RAND_424 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_166 = _RAND_424[21:0];
  _RAND_425 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_167 = _RAND_425[21:0];
  _RAND_426 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_168 = _RAND_426[21:0];
  _RAND_427 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_169 = _RAND_427[21:0];
  _RAND_428 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_170 = _RAND_428[21:0];
  _RAND_429 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_171 = _RAND_429[21:0];
  _RAND_430 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_172 = _RAND_430[21:0];
  _RAND_431 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_173 = _RAND_431[21:0];
  _RAND_432 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_174 = _RAND_432[21:0];
  _RAND_433 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_175 = _RAND_433[21:0];
  _RAND_434 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_176 = _RAND_434[21:0];
  _RAND_435 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_177 = _RAND_435[21:0];
  _RAND_436 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_178 = _RAND_436[21:0];
  _RAND_437 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_179 = _RAND_437[21:0];
  _RAND_438 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_180 = _RAND_438[21:0];
  _RAND_439 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_181 = _RAND_439[21:0];
  _RAND_440 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_182 = _RAND_440[21:0];
  _RAND_441 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_183 = _RAND_441[21:0];
  _RAND_442 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_184 = _RAND_442[21:0];
  _RAND_443 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_185 = _RAND_443[21:0];
  _RAND_444 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_186 = _RAND_444[21:0];
  _RAND_445 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_187 = _RAND_445[21:0];
  _RAND_446 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_188 = _RAND_446[21:0];
  _RAND_447 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_189 = _RAND_447[21:0];
  _RAND_448 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_190 = _RAND_448[21:0];
  _RAND_449 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_191 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_192 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_193 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_194 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_195 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_196 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_197 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_198 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_199 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_200 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_201 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_202 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_203 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_204 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_205 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_206 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_207 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_208 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_209 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_210 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_211 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_212 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_213 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_214 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_215 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_216 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_217 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_218 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_219 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_220 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_221 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_222 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_223 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_224 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_225 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_226 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_227 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_228 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_229 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_230 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_231 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_232 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_233 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_234 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_235 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_236 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_237 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_238 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_239 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_240 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_241 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_242 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_243 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_244 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_245 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_246 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_247 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_248 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_249 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_250 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_251 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_252 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_253 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_254 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_255 = _RAND_513[21:0];
  _RAND_514 = {1{`RANDOM}};
  fghr = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_0 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_1 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_2 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_3 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_4 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_5 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_6 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_7 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_8 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_9 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_10 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_11 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_12 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_13 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_14 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_15 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_16 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_17 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_18 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_19 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_20 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_21 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_22 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_23 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_24 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_25 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_26 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_27 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_28 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_29 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_30 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_31 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_32 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_33 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_34 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_35 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_36 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_37 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_38 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_39 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_40 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_41 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_42 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_43 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_44 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_45 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_46 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_47 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_48 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_49 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_50 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_51 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_52 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_53 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_54 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_55 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_56 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_57 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_58 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_59 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_60 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_61 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_62 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_63 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_64 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_65 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_66 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_67 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_68 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_69 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_70 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_71 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_72 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_73 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_74 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_75 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_76 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_77 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_78 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_79 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_80 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_81 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_82 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_83 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_84 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_85 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_86 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_87 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_88 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_89 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_90 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_91 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_92 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_93 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_94 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_95 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_96 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_97 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_98 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_99 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_100 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_101 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_102 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_103 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_104 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_105 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_106 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_107 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_108 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_109 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_110 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_111 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_112 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_113 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_114 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_115 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_116 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_117 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_118 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_119 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_120 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_121 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_122 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_123 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_124 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_125 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_126 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_127 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_128 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_129 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_130 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_131 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_132 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_133 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_134 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_135 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_136 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_137 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_138 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_139 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_140 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_141 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_142 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_143 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_144 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_145 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_146 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_147 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_148 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_149 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_150 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_151 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_152 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_153 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_154 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_155 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_156 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_157 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_158 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_159 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_160 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_161 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_162 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_163 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_164 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_165 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_166 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_167 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_168 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_169 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_170 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_171 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_172 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_173 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_174 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_175 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_176 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_177 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_178 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_179 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_180 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_181 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_182 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_183 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_184 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_185 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_186 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_187 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_188 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_189 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_190 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_191 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_192 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_193 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_194 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_195 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_196 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_197 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_198 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_199 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_200 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_201 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_202 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_203 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_204 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_205 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_206 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_207 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_208 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_209 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_210 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_211 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_212 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_213 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_214 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_215 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_216 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_217 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_218 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_219 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_220 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_221 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_222 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_223 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_224 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_225 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_226 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_227 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_228 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_229 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_230 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_231 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_232 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_233 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_234 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_235 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_236 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_237 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_238 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_239 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_240 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_241 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_242 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_243 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_244 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_245 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_246 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_247 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_248 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_249 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_250 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_251 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_252 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_253 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_254 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_255 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_0 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_1 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_2 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_3 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_4 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_5 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_6 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_7 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_8 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_9 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_10 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_11 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_12 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_13 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_14 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_15 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_16 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_17 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_18 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_19 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_20 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_21 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_22 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_23 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_24 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_25 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_26 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_27 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_28 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_29 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_30 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_31 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_32 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_33 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_34 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_35 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_36 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_37 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_38 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_39 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_40 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_41 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_42 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_43 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_44 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_45 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_46 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_47 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_48 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_49 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_50 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_51 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_52 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_53 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_54 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_55 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_56 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_57 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_58 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_59 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_60 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_61 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_62 = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_63 = _RAND_834[1:0];
  _RAND_835 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_64 = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_65 = _RAND_836[1:0];
  _RAND_837 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_66 = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_67 = _RAND_838[1:0];
  _RAND_839 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_68 = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_69 = _RAND_840[1:0];
  _RAND_841 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_70 = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_71 = _RAND_842[1:0];
  _RAND_843 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_72 = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_73 = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_74 = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_75 = _RAND_846[1:0];
  _RAND_847 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_76 = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_77 = _RAND_848[1:0];
  _RAND_849 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_78 = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_79 = _RAND_850[1:0];
  _RAND_851 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_80 = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_81 = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_82 = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_83 = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_84 = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_85 = _RAND_856[1:0];
  _RAND_857 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_86 = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_87 = _RAND_858[1:0];
  _RAND_859 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_88 = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_89 = _RAND_860[1:0];
  _RAND_861 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_90 = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_91 = _RAND_862[1:0];
  _RAND_863 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_92 = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_93 = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_94 = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_95 = _RAND_866[1:0];
  _RAND_867 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_96 = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_97 = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_98 = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_99 = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_100 = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_101 = _RAND_872[1:0];
  _RAND_873 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_102 = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_103 = _RAND_874[1:0];
  _RAND_875 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_104 = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_105 = _RAND_876[1:0];
  _RAND_877 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_106 = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_107 = _RAND_878[1:0];
  _RAND_879 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_108 = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_109 = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_110 = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_111 = _RAND_882[1:0];
  _RAND_883 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_112 = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_113 = _RAND_884[1:0];
  _RAND_885 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_114 = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_115 = _RAND_886[1:0];
  _RAND_887 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_116 = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_117 = _RAND_888[1:0];
  _RAND_889 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_118 = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_119 = _RAND_890[1:0];
  _RAND_891 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_120 = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_121 = _RAND_892[1:0];
  _RAND_893 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_122 = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_123 = _RAND_894[1:0];
  _RAND_895 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_124 = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_125 = _RAND_896[1:0];
  _RAND_897 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_126 = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_127 = _RAND_898[1:0];
  _RAND_899 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_128 = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_129 = _RAND_900[1:0];
  _RAND_901 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_130 = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_131 = _RAND_902[1:0];
  _RAND_903 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_132 = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_133 = _RAND_904[1:0];
  _RAND_905 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_134 = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_135 = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_136 = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_137 = _RAND_908[1:0];
  _RAND_909 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_138 = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_139 = _RAND_910[1:0];
  _RAND_911 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_140 = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_141 = _RAND_912[1:0];
  _RAND_913 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_142 = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_143 = _RAND_914[1:0];
  _RAND_915 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_144 = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_145 = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_146 = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_147 = _RAND_918[1:0];
  _RAND_919 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_148 = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_149 = _RAND_920[1:0];
  _RAND_921 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_150 = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_151 = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_152 = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_153 = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_154 = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_155 = _RAND_926[1:0];
  _RAND_927 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_156 = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_157 = _RAND_928[1:0];
  _RAND_929 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_158 = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_159 = _RAND_930[1:0];
  _RAND_931 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_160 = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_161 = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_162 = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_163 = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_164 = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_165 = _RAND_936[1:0];
  _RAND_937 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_166 = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_167 = _RAND_938[1:0];
  _RAND_939 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_168 = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_169 = _RAND_940[1:0];
  _RAND_941 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_170 = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_171 = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_172 = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_173 = _RAND_944[1:0];
  _RAND_945 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_174 = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_175 = _RAND_946[1:0];
  _RAND_947 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_176 = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_177 = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_178 = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_179 = _RAND_950[1:0];
  _RAND_951 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_180 = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_181 = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_182 = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_183 = _RAND_954[1:0];
  _RAND_955 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_184 = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_185 = _RAND_956[1:0];
  _RAND_957 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_186 = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_187 = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_188 = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_189 = _RAND_960[1:0];
  _RAND_961 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_190 = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_191 = _RAND_962[1:0];
  _RAND_963 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_192 = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_193 = _RAND_964[1:0];
  _RAND_965 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_194 = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_195 = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_196 = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_197 = _RAND_968[1:0];
  _RAND_969 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_198 = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_199 = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_200 = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_201 = _RAND_972[1:0];
  _RAND_973 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_202 = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_203 = _RAND_974[1:0];
  _RAND_975 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_204 = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_205 = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_206 = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_207 = _RAND_978[1:0];
  _RAND_979 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_208 = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_209 = _RAND_980[1:0];
  _RAND_981 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_210 = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_211 = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_212 = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_213 = _RAND_984[1:0];
  _RAND_985 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_214 = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_215 = _RAND_986[1:0];
  _RAND_987 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_216 = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_217 = _RAND_988[1:0];
  _RAND_989 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_218 = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_219 = _RAND_990[1:0];
  _RAND_991 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_220 = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_221 = _RAND_992[1:0];
  _RAND_993 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_222 = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_223 = _RAND_994[1:0];
  _RAND_995 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_224 = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_225 = _RAND_996[1:0];
  _RAND_997 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_226 = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_227 = _RAND_998[1:0];
  _RAND_999 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_228 = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_229 = _RAND_1000[1:0];
  _RAND_1001 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_230 = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_231 = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_232 = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_233 = _RAND_1004[1:0];
  _RAND_1005 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_234 = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_235 = _RAND_1006[1:0];
  _RAND_1007 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_236 = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_237 = _RAND_1008[1:0];
  _RAND_1009 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_238 = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_239 = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_240 = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_241 = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_242 = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_243 = _RAND_1014[1:0];
  _RAND_1015 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_244 = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_245 = _RAND_1016[1:0];
  _RAND_1017 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_246 = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_247 = _RAND_1018[1:0];
  _RAND_1019 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_248 = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_249 = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_250 = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_251 = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_252 = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_253 = _RAND_1024[1:0];
  _RAND_1025 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_254 = _RAND_1025[1:0];
  _RAND_1026 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_255 = _RAND_1026[1:0];
  _RAND_1027 = {1{`RANDOM}};
  exu_mp_way_f = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  exu_flush_final_d1 = _RAND_1028[0:0];
  _RAND_1029 = {8{`RANDOM}};
  btb_lru_b0_f = _RAND_1029[255:0];
  _RAND_1030 = {1{`RANDOM}};
  ifc_fetch_adder_prior = _RAND_1030[30:0];
  _RAND_1031 = {1{`RANDOM}};
  rets_out_0 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  rets_out_1 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  rets_out_2 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  rets_out_3 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  rets_out_4 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  rets_out_5 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  rets_out_6 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  rets_out_7 = _RAND_1038[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    leak_one_f_d1 = 1'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_255 = 22'h0;
  end
  if (reset) begin
    dec_tlu_way_wb_f = 1'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_255 = 22'h0;
  end
  if (reset) begin
    fghr = 8'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_255 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_255 = 2'h0;
  end
  if (reset) begin
    exu_mp_way_f = 1'h0;
  end
  if (reset) begin
    exu_flush_final_d1 = 1'h0;
  end
  if (reset) begin
    btb_lru_b0_f = 256'h0;
  end
  if (reset) begin
    ifc_fetch_adder_prior = 31'h0;
  end
  if (reset) begin
    rets_out_0 = 32'h0;
  end
  if (reset) begin
    rets_out_1 = 32'h0;
  end
  if (reset) begin
    rets_out_2 = 32'h0;
  end
  if (reset) begin
    rets_out_3 = 32'h0;
  end
  if (reset) begin
    rets_out_4 = 32'h0;
  end
  if (reset) begin
    rets_out_5 = 32'h0;
  end
  if (reset) begin
    rets_out_6 = 32'h0;
  end
  if (reset) begin
    rets_out_7 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      leak_one_f_d1 <= 1'h0;
    end else begin
      leak_one_f_d1 <= _T_40 | _T_41;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_0 <= 22'h0;
    end else if (_T_573) begin
      btb_bank0_rd_data_way0_out_0 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_1 <= 22'h0;
    end else if (_T_576) begin
      btb_bank0_rd_data_way0_out_1 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_2 <= 22'h0;
    end else if (_T_579) begin
      btb_bank0_rd_data_way0_out_2 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_3 <= 22'h0;
    end else if (_T_582) begin
      btb_bank0_rd_data_way0_out_3 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_4 <= 22'h0;
    end else if (_T_585) begin
      btb_bank0_rd_data_way0_out_4 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_5 <= 22'h0;
    end else if (_T_588) begin
      btb_bank0_rd_data_way0_out_5 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_6 <= 22'h0;
    end else if (_T_591) begin
      btb_bank0_rd_data_way0_out_6 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_7 <= 22'h0;
    end else if (_T_594) begin
      btb_bank0_rd_data_way0_out_7 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_8 <= 22'h0;
    end else if (_T_597) begin
      btb_bank0_rd_data_way0_out_8 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_9 <= 22'h0;
    end else if (_T_600) begin
      btb_bank0_rd_data_way0_out_9 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_10 <= 22'h0;
    end else if (_T_603) begin
      btb_bank0_rd_data_way0_out_10 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_11 <= 22'h0;
    end else if (_T_606) begin
      btb_bank0_rd_data_way0_out_11 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_12 <= 22'h0;
    end else if (_T_609) begin
      btb_bank0_rd_data_way0_out_12 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_13 <= 22'h0;
    end else if (_T_612) begin
      btb_bank0_rd_data_way0_out_13 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_14 <= 22'h0;
    end else if (_T_615) begin
      btb_bank0_rd_data_way0_out_14 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_15 <= 22'h0;
    end else if (_T_618) begin
      btb_bank0_rd_data_way0_out_15 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_16 <= 22'h0;
    end else if (_T_621) begin
      btb_bank0_rd_data_way0_out_16 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_17 <= 22'h0;
    end else if (_T_624) begin
      btb_bank0_rd_data_way0_out_17 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_18 <= 22'h0;
    end else if (_T_627) begin
      btb_bank0_rd_data_way0_out_18 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_19 <= 22'h0;
    end else if (_T_630) begin
      btb_bank0_rd_data_way0_out_19 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_20 <= 22'h0;
    end else if (_T_633) begin
      btb_bank0_rd_data_way0_out_20 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_21 <= 22'h0;
    end else if (_T_636) begin
      btb_bank0_rd_data_way0_out_21 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_22 <= 22'h0;
    end else if (_T_639) begin
      btb_bank0_rd_data_way0_out_22 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_23 <= 22'h0;
    end else if (_T_642) begin
      btb_bank0_rd_data_way0_out_23 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_24 <= 22'h0;
    end else if (_T_645) begin
      btb_bank0_rd_data_way0_out_24 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_25 <= 22'h0;
    end else if (_T_648) begin
      btb_bank0_rd_data_way0_out_25 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_26 <= 22'h0;
    end else if (_T_651) begin
      btb_bank0_rd_data_way0_out_26 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_27 <= 22'h0;
    end else if (_T_654) begin
      btb_bank0_rd_data_way0_out_27 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_28 <= 22'h0;
    end else if (_T_657) begin
      btb_bank0_rd_data_way0_out_28 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_29 <= 22'h0;
    end else if (_T_660) begin
      btb_bank0_rd_data_way0_out_29 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_30 <= 22'h0;
    end else if (_T_663) begin
      btb_bank0_rd_data_way0_out_30 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_31 <= 22'h0;
    end else if (_T_666) begin
      btb_bank0_rd_data_way0_out_31 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_32 <= 22'h0;
    end else if (_T_669) begin
      btb_bank0_rd_data_way0_out_32 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_33 <= 22'h0;
    end else if (_T_672) begin
      btb_bank0_rd_data_way0_out_33 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_34 <= 22'h0;
    end else if (_T_675) begin
      btb_bank0_rd_data_way0_out_34 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_35 <= 22'h0;
    end else if (_T_678) begin
      btb_bank0_rd_data_way0_out_35 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_36 <= 22'h0;
    end else if (_T_681) begin
      btb_bank0_rd_data_way0_out_36 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_37 <= 22'h0;
    end else if (_T_684) begin
      btb_bank0_rd_data_way0_out_37 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_38 <= 22'h0;
    end else if (_T_687) begin
      btb_bank0_rd_data_way0_out_38 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_39 <= 22'h0;
    end else if (_T_690) begin
      btb_bank0_rd_data_way0_out_39 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_40 <= 22'h0;
    end else if (_T_693) begin
      btb_bank0_rd_data_way0_out_40 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_41 <= 22'h0;
    end else if (_T_696) begin
      btb_bank0_rd_data_way0_out_41 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_42 <= 22'h0;
    end else if (_T_699) begin
      btb_bank0_rd_data_way0_out_42 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_43 <= 22'h0;
    end else if (_T_702) begin
      btb_bank0_rd_data_way0_out_43 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_44 <= 22'h0;
    end else if (_T_705) begin
      btb_bank0_rd_data_way0_out_44 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_45 <= 22'h0;
    end else if (_T_708) begin
      btb_bank0_rd_data_way0_out_45 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_46 <= 22'h0;
    end else if (_T_711) begin
      btb_bank0_rd_data_way0_out_46 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_47 <= 22'h0;
    end else if (_T_714) begin
      btb_bank0_rd_data_way0_out_47 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_48 <= 22'h0;
    end else if (_T_717) begin
      btb_bank0_rd_data_way0_out_48 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_49 <= 22'h0;
    end else if (_T_720) begin
      btb_bank0_rd_data_way0_out_49 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_50 <= 22'h0;
    end else if (_T_723) begin
      btb_bank0_rd_data_way0_out_50 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_51 <= 22'h0;
    end else if (_T_726) begin
      btb_bank0_rd_data_way0_out_51 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_52 <= 22'h0;
    end else if (_T_729) begin
      btb_bank0_rd_data_way0_out_52 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_53 <= 22'h0;
    end else if (_T_732) begin
      btb_bank0_rd_data_way0_out_53 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_54 <= 22'h0;
    end else if (_T_735) begin
      btb_bank0_rd_data_way0_out_54 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_55 <= 22'h0;
    end else if (_T_738) begin
      btb_bank0_rd_data_way0_out_55 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_56 <= 22'h0;
    end else if (_T_741) begin
      btb_bank0_rd_data_way0_out_56 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_57 <= 22'h0;
    end else if (_T_744) begin
      btb_bank0_rd_data_way0_out_57 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_58 <= 22'h0;
    end else if (_T_747) begin
      btb_bank0_rd_data_way0_out_58 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_59 <= 22'h0;
    end else if (_T_750) begin
      btb_bank0_rd_data_way0_out_59 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_60 <= 22'h0;
    end else if (_T_753) begin
      btb_bank0_rd_data_way0_out_60 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_61 <= 22'h0;
    end else if (_T_756) begin
      btb_bank0_rd_data_way0_out_61 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_62 <= 22'h0;
    end else if (_T_759) begin
      btb_bank0_rd_data_way0_out_62 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_63 <= 22'h0;
    end else if (_T_762) begin
      btb_bank0_rd_data_way0_out_63 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_64 <= 22'h0;
    end else if (_T_765) begin
      btb_bank0_rd_data_way0_out_64 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_65 <= 22'h0;
    end else if (_T_768) begin
      btb_bank0_rd_data_way0_out_65 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_66 <= 22'h0;
    end else if (_T_771) begin
      btb_bank0_rd_data_way0_out_66 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_67 <= 22'h0;
    end else if (_T_774) begin
      btb_bank0_rd_data_way0_out_67 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_68 <= 22'h0;
    end else if (_T_777) begin
      btb_bank0_rd_data_way0_out_68 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_69 <= 22'h0;
    end else if (_T_780) begin
      btb_bank0_rd_data_way0_out_69 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_70 <= 22'h0;
    end else if (_T_783) begin
      btb_bank0_rd_data_way0_out_70 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_71 <= 22'h0;
    end else if (_T_786) begin
      btb_bank0_rd_data_way0_out_71 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_72 <= 22'h0;
    end else if (_T_789) begin
      btb_bank0_rd_data_way0_out_72 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_73 <= 22'h0;
    end else if (_T_792) begin
      btb_bank0_rd_data_way0_out_73 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_74 <= 22'h0;
    end else if (_T_795) begin
      btb_bank0_rd_data_way0_out_74 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_75 <= 22'h0;
    end else if (_T_798) begin
      btb_bank0_rd_data_way0_out_75 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_76 <= 22'h0;
    end else if (_T_801) begin
      btb_bank0_rd_data_way0_out_76 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_77 <= 22'h0;
    end else if (_T_804) begin
      btb_bank0_rd_data_way0_out_77 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_78 <= 22'h0;
    end else if (_T_807) begin
      btb_bank0_rd_data_way0_out_78 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_79 <= 22'h0;
    end else if (_T_810) begin
      btb_bank0_rd_data_way0_out_79 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_80 <= 22'h0;
    end else if (_T_813) begin
      btb_bank0_rd_data_way0_out_80 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_81 <= 22'h0;
    end else if (_T_816) begin
      btb_bank0_rd_data_way0_out_81 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_82 <= 22'h0;
    end else if (_T_819) begin
      btb_bank0_rd_data_way0_out_82 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_83 <= 22'h0;
    end else if (_T_822) begin
      btb_bank0_rd_data_way0_out_83 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_84 <= 22'h0;
    end else if (_T_825) begin
      btb_bank0_rd_data_way0_out_84 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_85 <= 22'h0;
    end else if (_T_828) begin
      btb_bank0_rd_data_way0_out_85 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_86 <= 22'h0;
    end else if (_T_831) begin
      btb_bank0_rd_data_way0_out_86 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_87 <= 22'h0;
    end else if (_T_834) begin
      btb_bank0_rd_data_way0_out_87 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_88 <= 22'h0;
    end else if (_T_837) begin
      btb_bank0_rd_data_way0_out_88 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_89 <= 22'h0;
    end else if (_T_840) begin
      btb_bank0_rd_data_way0_out_89 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_90 <= 22'h0;
    end else if (_T_843) begin
      btb_bank0_rd_data_way0_out_90 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_91 <= 22'h0;
    end else if (_T_846) begin
      btb_bank0_rd_data_way0_out_91 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_92 <= 22'h0;
    end else if (_T_849) begin
      btb_bank0_rd_data_way0_out_92 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_93 <= 22'h0;
    end else if (_T_852) begin
      btb_bank0_rd_data_way0_out_93 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_94 <= 22'h0;
    end else if (_T_855) begin
      btb_bank0_rd_data_way0_out_94 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_95 <= 22'h0;
    end else if (_T_858) begin
      btb_bank0_rd_data_way0_out_95 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_96 <= 22'h0;
    end else if (_T_861) begin
      btb_bank0_rd_data_way0_out_96 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_97 <= 22'h0;
    end else if (_T_864) begin
      btb_bank0_rd_data_way0_out_97 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_98 <= 22'h0;
    end else if (_T_867) begin
      btb_bank0_rd_data_way0_out_98 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_99 <= 22'h0;
    end else if (_T_870) begin
      btb_bank0_rd_data_way0_out_99 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_100 <= 22'h0;
    end else if (_T_873) begin
      btb_bank0_rd_data_way0_out_100 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_101 <= 22'h0;
    end else if (_T_876) begin
      btb_bank0_rd_data_way0_out_101 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_102 <= 22'h0;
    end else if (_T_879) begin
      btb_bank0_rd_data_way0_out_102 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_103 <= 22'h0;
    end else if (_T_882) begin
      btb_bank0_rd_data_way0_out_103 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_104 <= 22'h0;
    end else if (_T_885) begin
      btb_bank0_rd_data_way0_out_104 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_105 <= 22'h0;
    end else if (_T_888) begin
      btb_bank0_rd_data_way0_out_105 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_106 <= 22'h0;
    end else if (_T_891) begin
      btb_bank0_rd_data_way0_out_106 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_107 <= 22'h0;
    end else if (_T_894) begin
      btb_bank0_rd_data_way0_out_107 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_108 <= 22'h0;
    end else if (_T_897) begin
      btb_bank0_rd_data_way0_out_108 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_109 <= 22'h0;
    end else if (_T_900) begin
      btb_bank0_rd_data_way0_out_109 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_110 <= 22'h0;
    end else if (_T_903) begin
      btb_bank0_rd_data_way0_out_110 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_111 <= 22'h0;
    end else if (_T_906) begin
      btb_bank0_rd_data_way0_out_111 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_112 <= 22'h0;
    end else if (_T_909) begin
      btb_bank0_rd_data_way0_out_112 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_113 <= 22'h0;
    end else if (_T_912) begin
      btb_bank0_rd_data_way0_out_113 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_114 <= 22'h0;
    end else if (_T_915) begin
      btb_bank0_rd_data_way0_out_114 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_115 <= 22'h0;
    end else if (_T_918) begin
      btb_bank0_rd_data_way0_out_115 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_116 <= 22'h0;
    end else if (_T_921) begin
      btb_bank0_rd_data_way0_out_116 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_117 <= 22'h0;
    end else if (_T_924) begin
      btb_bank0_rd_data_way0_out_117 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_118 <= 22'h0;
    end else if (_T_927) begin
      btb_bank0_rd_data_way0_out_118 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_119 <= 22'h0;
    end else if (_T_930) begin
      btb_bank0_rd_data_way0_out_119 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_120 <= 22'h0;
    end else if (_T_933) begin
      btb_bank0_rd_data_way0_out_120 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_121 <= 22'h0;
    end else if (_T_936) begin
      btb_bank0_rd_data_way0_out_121 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_122 <= 22'h0;
    end else if (_T_939) begin
      btb_bank0_rd_data_way0_out_122 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_123 <= 22'h0;
    end else if (_T_942) begin
      btb_bank0_rd_data_way0_out_123 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_124 <= 22'h0;
    end else if (_T_945) begin
      btb_bank0_rd_data_way0_out_124 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_125 <= 22'h0;
    end else if (_T_948) begin
      btb_bank0_rd_data_way0_out_125 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_126 <= 22'h0;
    end else if (_T_951) begin
      btb_bank0_rd_data_way0_out_126 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_127 <= 22'h0;
    end else if (_T_954) begin
      btb_bank0_rd_data_way0_out_127 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_128 <= 22'h0;
    end else if (_T_957) begin
      btb_bank0_rd_data_way0_out_128 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_129 <= 22'h0;
    end else if (_T_960) begin
      btb_bank0_rd_data_way0_out_129 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_130 <= 22'h0;
    end else if (_T_963) begin
      btb_bank0_rd_data_way0_out_130 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_131 <= 22'h0;
    end else if (_T_966) begin
      btb_bank0_rd_data_way0_out_131 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_132 <= 22'h0;
    end else if (_T_969) begin
      btb_bank0_rd_data_way0_out_132 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_133 <= 22'h0;
    end else if (_T_972) begin
      btb_bank0_rd_data_way0_out_133 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_134 <= 22'h0;
    end else if (_T_975) begin
      btb_bank0_rd_data_way0_out_134 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_135 <= 22'h0;
    end else if (_T_978) begin
      btb_bank0_rd_data_way0_out_135 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_136 <= 22'h0;
    end else if (_T_981) begin
      btb_bank0_rd_data_way0_out_136 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_137 <= 22'h0;
    end else if (_T_984) begin
      btb_bank0_rd_data_way0_out_137 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_138 <= 22'h0;
    end else if (_T_987) begin
      btb_bank0_rd_data_way0_out_138 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_139 <= 22'h0;
    end else if (_T_990) begin
      btb_bank0_rd_data_way0_out_139 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_140 <= 22'h0;
    end else if (_T_993) begin
      btb_bank0_rd_data_way0_out_140 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_141 <= 22'h0;
    end else if (_T_996) begin
      btb_bank0_rd_data_way0_out_141 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_142 <= 22'h0;
    end else if (_T_999) begin
      btb_bank0_rd_data_way0_out_142 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_143 <= 22'h0;
    end else if (_T_1002) begin
      btb_bank0_rd_data_way0_out_143 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_144 <= 22'h0;
    end else if (_T_1005) begin
      btb_bank0_rd_data_way0_out_144 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_145 <= 22'h0;
    end else if (_T_1008) begin
      btb_bank0_rd_data_way0_out_145 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_146 <= 22'h0;
    end else if (_T_1011) begin
      btb_bank0_rd_data_way0_out_146 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_147 <= 22'h0;
    end else if (_T_1014) begin
      btb_bank0_rd_data_way0_out_147 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_148 <= 22'h0;
    end else if (_T_1017) begin
      btb_bank0_rd_data_way0_out_148 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_149 <= 22'h0;
    end else if (_T_1020) begin
      btb_bank0_rd_data_way0_out_149 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_150 <= 22'h0;
    end else if (_T_1023) begin
      btb_bank0_rd_data_way0_out_150 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_151 <= 22'h0;
    end else if (_T_1026) begin
      btb_bank0_rd_data_way0_out_151 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_152 <= 22'h0;
    end else if (_T_1029) begin
      btb_bank0_rd_data_way0_out_152 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_153 <= 22'h0;
    end else if (_T_1032) begin
      btb_bank0_rd_data_way0_out_153 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_154 <= 22'h0;
    end else if (_T_1035) begin
      btb_bank0_rd_data_way0_out_154 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_155 <= 22'h0;
    end else if (_T_1038) begin
      btb_bank0_rd_data_way0_out_155 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_156 <= 22'h0;
    end else if (_T_1041) begin
      btb_bank0_rd_data_way0_out_156 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_157 <= 22'h0;
    end else if (_T_1044) begin
      btb_bank0_rd_data_way0_out_157 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_158 <= 22'h0;
    end else if (_T_1047) begin
      btb_bank0_rd_data_way0_out_158 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_159 <= 22'h0;
    end else if (_T_1050) begin
      btb_bank0_rd_data_way0_out_159 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_160 <= 22'h0;
    end else if (_T_1053) begin
      btb_bank0_rd_data_way0_out_160 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_161 <= 22'h0;
    end else if (_T_1056) begin
      btb_bank0_rd_data_way0_out_161 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_162 <= 22'h0;
    end else if (_T_1059) begin
      btb_bank0_rd_data_way0_out_162 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_163 <= 22'h0;
    end else if (_T_1062) begin
      btb_bank0_rd_data_way0_out_163 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_164 <= 22'h0;
    end else if (_T_1065) begin
      btb_bank0_rd_data_way0_out_164 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_165 <= 22'h0;
    end else if (_T_1068) begin
      btb_bank0_rd_data_way0_out_165 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_166 <= 22'h0;
    end else if (_T_1071) begin
      btb_bank0_rd_data_way0_out_166 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_167 <= 22'h0;
    end else if (_T_1074) begin
      btb_bank0_rd_data_way0_out_167 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_168 <= 22'h0;
    end else if (_T_1077) begin
      btb_bank0_rd_data_way0_out_168 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_169 <= 22'h0;
    end else if (_T_1080) begin
      btb_bank0_rd_data_way0_out_169 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_170 <= 22'h0;
    end else if (_T_1083) begin
      btb_bank0_rd_data_way0_out_170 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_171 <= 22'h0;
    end else if (_T_1086) begin
      btb_bank0_rd_data_way0_out_171 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_172 <= 22'h0;
    end else if (_T_1089) begin
      btb_bank0_rd_data_way0_out_172 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_173 <= 22'h0;
    end else if (_T_1092) begin
      btb_bank0_rd_data_way0_out_173 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_174 <= 22'h0;
    end else if (_T_1095) begin
      btb_bank0_rd_data_way0_out_174 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_175 <= 22'h0;
    end else if (_T_1098) begin
      btb_bank0_rd_data_way0_out_175 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_176 <= 22'h0;
    end else if (_T_1101) begin
      btb_bank0_rd_data_way0_out_176 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_177 <= 22'h0;
    end else if (_T_1104) begin
      btb_bank0_rd_data_way0_out_177 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_178 <= 22'h0;
    end else if (_T_1107) begin
      btb_bank0_rd_data_way0_out_178 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_179 <= 22'h0;
    end else if (_T_1110) begin
      btb_bank0_rd_data_way0_out_179 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_180 <= 22'h0;
    end else if (_T_1113) begin
      btb_bank0_rd_data_way0_out_180 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_181 <= 22'h0;
    end else if (_T_1116) begin
      btb_bank0_rd_data_way0_out_181 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_182 <= 22'h0;
    end else if (_T_1119) begin
      btb_bank0_rd_data_way0_out_182 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_183 <= 22'h0;
    end else if (_T_1122) begin
      btb_bank0_rd_data_way0_out_183 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_184 <= 22'h0;
    end else if (_T_1125) begin
      btb_bank0_rd_data_way0_out_184 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_185 <= 22'h0;
    end else if (_T_1128) begin
      btb_bank0_rd_data_way0_out_185 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_186 <= 22'h0;
    end else if (_T_1131) begin
      btb_bank0_rd_data_way0_out_186 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_187 <= 22'h0;
    end else if (_T_1134) begin
      btb_bank0_rd_data_way0_out_187 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_188 <= 22'h0;
    end else if (_T_1137) begin
      btb_bank0_rd_data_way0_out_188 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_189 <= 22'h0;
    end else if (_T_1140) begin
      btb_bank0_rd_data_way0_out_189 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_190 <= 22'h0;
    end else if (_T_1143) begin
      btb_bank0_rd_data_way0_out_190 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_191 <= 22'h0;
    end else if (_T_1146) begin
      btb_bank0_rd_data_way0_out_191 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_192 <= 22'h0;
    end else if (_T_1149) begin
      btb_bank0_rd_data_way0_out_192 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_193 <= 22'h0;
    end else if (_T_1152) begin
      btb_bank0_rd_data_way0_out_193 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_194 <= 22'h0;
    end else if (_T_1155) begin
      btb_bank0_rd_data_way0_out_194 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_195 <= 22'h0;
    end else if (_T_1158) begin
      btb_bank0_rd_data_way0_out_195 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_196 <= 22'h0;
    end else if (_T_1161) begin
      btb_bank0_rd_data_way0_out_196 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_197 <= 22'h0;
    end else if (_T_1164) begin
      btb_bank0_rd_data_way0_out_197 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_198 <= 22'h0;
    end else if (_T_1167) begin
      btb_bank0_rd_data_way0_out_198 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_199 <= 22'h0;
    end else if (_T_1170) begin
      btb_bank0_rd_data_way0_out_199 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_200 <= 22'h0;
    end else if (_T_1173) begin
      btb_bank0_rd_data_way0_out_200 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_201 <= 22'h0;
    end else if (_T_1176) begin
      btb_bank0_rd_data_way0_out_201 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_202 <= 22'h0;
    end else if (_T_1179) begin
      btb_bank0_rd_data_way0_out_202 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_203 <= 22'h0;
    end else if (_T_1182) begin
      btb_bank0_rd_data_way0_out_203 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_204 <= 22'h0;
    end else if (_T_1185) begin
      btb_bank0_rd_data_way0_out_204 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_205 <= 22'h0;
    end else if (_T_1188) begin
      btb_bank0_rd_data_way0_out_205 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_206 <= 22'h0;
    end else if (_T_1191) begin
      btb_bank0_rd_data_way0_out_206 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_207 <= 22'h0;
    end else if (_T_1194) begin
      btb_bank0_rd_data_way0_out_207 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_208 <= 22'h0;
    end else if (_T_1197) begin
      btb_bank0_rd_data_way0_out_208 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_209 <= 22'h0;
    end else if (_T_1200) begin
      btb_bank0_rd_data_way0_out_209 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_210 <= 22'h0;
    end else if (_T_1203) begin
      btb_bank0_rd_data_way0_out_210 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_211 <= 22'h0;
    end else if (_T_1206) begin
      btb_bank0_rd_data_way0_out_211 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_212 <= 22'h0;
    end else if (_T_1209) begin
      btb_bank0_rd_data_way0_out_212 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_213 <= 22'h0;
    end else if (_T_1212) begin
      btb_bank0_rd_data_way0_out_213 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_214 <= 22'h0;
    end else if (_T_1215) begin
      btb_bank0_rd_data_way0_out_214 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_215 <= 22'h0;
    end else if (_T_1218) begin
      btb_bank0_rd_data_way0_out_215 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_216 <= 22'h0;
    end else if (_T_1221) begin
      btb_bank0_rd_data_way0_out_216 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_217 <= 22'h0;
    end else if (_T_1224) begin
      btb_bank0_rd_data_way0_out_217 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_218 <= 22'h0;
    end else if (_T_1227) begin
      btb_bank0_rd_data_way0_out_218 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_219 <= 22'h0;
    end else if (_T_1230) begin
      btb_bank0_rd_data_way0_out_219 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_220 <= 22'h0;
    end else if (_T_1233) begin
      btb_bank0_rd_data_way0_out_220 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_221 <= 22'h0;
    end else if (_T_1236) begin
      btb_bank0_rd_data_way0_out_221 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_222 <= 22'h0;
    end else if (_T_1239) begin
      btb_bank0_rd_data_way0_out_222 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_223 <= 22'h0;
    end else if (_T_1242) begin
      btb_bank0_rd_data_way0_out_223 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_224 <= 22'h0;
    end else if (_T_1245) begin
      btb_bank0_rd_data_way0_out_224 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_225 <= 22'h0;
    end else if (_T_1248) begin
      btb_bank0_rd_data_way0_out_225 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_226 <= 22'h0;
    end else if (_T_1251) begin
      btb_bank0_rd_data_way0_out_226 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_227 <= 22'h0;
    end else if (_T_1254) begin
      btb_bank0_rd_data_way0_out_227 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_228 <= 22'h0;
    end else if (_T_1257) begin
      btb_bank0_rd_data_way0_out_228 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_229 <= 22'h0;
    end else if (_T_1260) begin
      btb_bank0_rd_data_way0_out_229 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_230 <= 22'h0;
    end else if (_T_1263) begin
      btb_bank0_rd_data_way0_out_230 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_231 <= 22'h0;
    end else if (_T_1266) begin
      btb_bank0_rd_data_way0_out_231 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_232 <= 22'h0;
    end else if (_T_1269) begin
      btb_bank0_rd_data_way0_out_232 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_233 <= 22'h0;
    end else if (_T_1272) begin
      btb_bank0_rd_data_way0_out_233 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_234 <= 22'h0;
    end else if (_T_1275) begin
      btb_bank0_rd_data_way0_out_234 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_235 <= 22'h0;
    end else if (_T_1278) begin
      btb_bank0_rd_data_way0_out_235 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_236 <= 22'h0;
    end else if (_T_1281) begin
      btb_bank0_rd_data_way0_out_236 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_237 <= 22'h0;
    end else if (_T_1284) begin
      btb_bank0_rd_data_way0_out_237 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_238 <= 22'h0;
    end else if (_T_1287) begin
      btb_bank0_rd_data_way0_out_238 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_239 <= 22'h0;
    end else if (_T_1290) begin
      btb_bank0_rd_data_way0_out_239 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_240 <= 22'h0;
    end else if (_T_1293) begin
      btb_bank0_rd_data_way0_out_240 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_241 <= 22'h0;
    end else if (_T_1296) begin
      btb_bank0_rd_data_way0_out_241 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_242 <= 22'h0;
    end else if (_T_1299) begin
      btb_bank0_rd_data_way0_out_242 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_243 <= 22'h0;
    end else if (_T_1302) begin
      btb_bank0_rd_data_way0_out_243 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_244 <= 22'h0;
    end else if (_T_1305) begin
      btb_bank0_rd_data_way0_out_244 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_245 <= 22'h0;
    end else if (_T_1308) begin
      btb_bank0_rd_data_way0_out_245 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_246 <= 22'h0;
    end else if (_T_1311) begin
      btb_bank0_rd_data_way0_out_246 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_247 <= 22'h0;
    end else if (_T_1314) begin
      btb_bank0_rd_data_way0_out_247 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_248 <= 22'h0;
    end else if (_T_1317) begin
      btb_bank0_rd_data_way0_out_248 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_249 <= 22'h0;
    end else if (_T_1320) begin
      btb_bank0_rd_data_way0_out_249 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_250 <= 22'h0;
    end else if (_T_1323) begin
      btb_bank0_rd_data_way0_out_250 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_251 <= 22'h0;
    end else if (_T_1326) begin
      btb_bank0_rd_data_way0_out_251 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_252 <= 22'h0;
    end else if (_T_1329) begin
      btb_bank0_rd_data_way0_out_252 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_253 <= 22'h0;
    end else if (_T_1332) begin
      btb_bank0_rd_data_way0_out_253 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_254 <= 22'h0;
    end else if (_T_1335) begin
      btb_bank0_rd_data_way0_out_254 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_255 <= 22'h0;
    end else if (_T_1338) begin
      btb_bank0_rd_data_way0_out_255 <= btb_wr_data;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      dec_tlu_way_wb_f <= 1'h0;
    end else begin
      dec_tlu_way_wb_f <= io_dec_tlu_br0_r_pkt_way;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_0 <= 22'h0;
    end else if (_T_1341) begin
      btb_bank0_rd_data_way1_out_0 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_1 <= 22'h0;
    end else if (_T_1344) begin
      btb_bank0_rd_data_way1_out_1 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_2 <= 22'h0;
    end else if (_T_1347) begin
      btb_bank0_rd_data_way1_out_2 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_3 <= 22'h0;
    end else if (_T_1350) begin
      btb_bank0_rd_data_way1_out_3 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_4 <= 22'h0;
    end else if (_T_1353) begin
      btb_bank0_rd_data_way1_out_4 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_5 <= 22'h0;
    end else if (_T_1356) begin
      btb_bank0_rd_data_way1_out_5 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_6 <= 22'h0;
    end else if (_T_1359) begin
      btb_bank0_rd_data_way1_out_6 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_7 <= 22'h0;
    end else if (_T_1362) begin
      btb_bank0_rd_data_way1_out_7 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_8 <= 22'h0;
    end else if (_T_1365) begin
      btb_bank0_rd_data_way1_out_8 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_9 <= 22'h0;
    end else if (_T_1368) begin
      btb_bank0_rd_data_way1_out_9 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_10 <= 22'h0;
    end else if (_T_1371) begin
      btb_bank0_rd_data_way1_out_10 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_11 <= 22'h0;
    end else if (_T_1374) begin
      btb_bank0_rd_data_way1_out_11 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_12 <= 22'h0;
    end else if (_T_1377) begin
      btb_bank0_rd_data_way1_out_12 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_13 <= 22'h0;
    end else if (_T_1380) begin
      btb_bank0_rd_data_way1_out_13 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_14 <= 22'h0;
    end else if (_T_1383) begin
      btb_bank0_rd_data_way1_out_14 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_15 <= 22'h0;
    end else if (_T_1386) begin
      btb_bank0_rd_data_way1_out_15 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_16 <= 22'h0;
    end else if (_T_1389) begin
      btb_bank0_rd_data_way1_out_16 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_17 <= 22'h0;
    end else if (_T_1392) begin
      btb_bank0_rd_data_way1_out_17 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_18 <= 22'h0;
    end else if (_T_1395) begin
      btb_bank0_rd_data_way1_out_18 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_19 <= 22'h0;
    end else if (_T_1398) begin
      btb_bank0_rd_data_way1_out_19 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_20 <= 22'h0;
    end else if (_T_1401) begin
      btb_bank0_rd_data_way1_out_20 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_21 <= 22'h0;
    end else if (_T_1404) begin
      btb_bank0_rd_data_way1_out_21 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_22 <= 22'h0;
    end else if (_T_1407) begin
      btb_bank0_rd_data_way1_out_22 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_23 <= 22'h0;
    end else if (_T_1410) begin
      btb_bank0_rd_data_way1_out_23 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_24 <= 22'h0;
    end else if (_T_1413) begin
      btb_bank0_rd_data_way1_out_24 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_25 <= 22'h0;
    end else if (_T_1416) begin
      btb_bank0_rd_data_way1_out_25 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_26 <= 22'h0;
    end else if (_T_1419) begin
      btb_bank0_rd_data_way1_out_26 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_27 <= 22'h0;
    end else if (_T_1422) begin
      btb_bank0_rd_data_way1_out_27 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_28 <= 22'h0;
    end else if (_T_1425) begin
      btb_bank0_rd_data_way1_out_28 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_29 <= 22'h0;
    end else if (_T_1428) begin
      btb_bank0_rd_data_way1_out_29 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_30 <= 22'h0;
    end else if (_T_1431) begin
      btb_bank0_rd_data_way1_out_30 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_31 <= 22'h0;
    end else if (_T_1434) begin
      btb_bank0_rd_data_way1_out_31 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_32 <= 22'h0;
    end else if (_T_1437) begin
      btb_bank0_rd_data_way1_out_32 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_33 <= 22'h0;
    end else if (_T_1440) begin
      btb_bank0_rd_data_way1_out_33 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_34 <= 22'h0;
    end else if (_T_1443) begin
      btb_bank0_rd_data_way1_out_34 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_35 <= 22'h0;
    end else if (_T_1446) begin
      btb_bank0_rd_data_way1_out_35 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_36 <= 22'h0;
    end else if (_T_1449) begin
      btb_bank0_rd_data_way1_out_36 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_37 <= 22'h0;
    end else if (_T_1452) begin
      btb_bank0_rd_data_way1_out_37 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_38 <= 22'h0;
    end else if (_T_1455) begin
      btb_bank0_rd_data_way1_out_38 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_39 <= 22'h0;
    end else if (_T_1458) begin
      btb_bank0_rd_data_way1_out_39 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_40 <= 22'h0;
    end else if (_T_1461) begin
      btb_bank0_rd_data_way1_out_40 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_41 <= 22'h0;
    end else if (_T_1464) begin
      btb_bank0_rd_data_way1_out_41 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_42 <= 22'h0;
    end else if (_T_1467) begin
      btb_bank0_rd_data_way1_out_42 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_43 <= 22'h0;
    end else if (_T_1470) begin
      btb_bank0_rd_data_way1_out_43 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_44 <= 22'h0;
    end else if (_T_1473) begin
      btb_bank0_rd_data_way1_out_44 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_45 <= 22'h0;
    end else if (_T_1476) begin
      btb_bank0_rd_data_way1_out_45 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_46 <= 22'h0;
    end else if (_T_1479) begin
      btb_bank0_rd_data_way1_out_46 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_47 <= 22'h0;
    end else if (_T_1482) begin
      btb_bank0_rd_data_way1_out_47 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_48 <= 22'h0;
    end else if (_T_1485) begin
      btb_bank0_rd_data_way1_out_48 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_49 <= 22'h0;
    end else if (_T_1488) begin
      btb_bank0_rd_data_way1_out_49 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_50 <= 22'h0;
    end else if (_T_1491) begin
      btb_bank0_rd_data_way1_out_50 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_51 <= 22'h0;
    end else if (_T_1494) begin
      btb_bank0_rd_data_way1_out_51 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_52 <= 22'h0;
    end else if (_T_1497) begin
      btb_bank0_rd_data_way1_out_52 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_53 <= 22'h0;
    end else if (_T_1500) begin
      btb_bank0_rd_data_way1_out_53 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_54 <= 22'h0;
    end else if (_T_1503) begin
      btb_bank0_rd_data_way1_out_54 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_55 <= 22'h0;
    end else if (_T_1506) begin
      btb_bank0_rd_data_way1_out_55 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_56 <= 22'h0;
    end else if (_T_1509) begin
      btb_bank0_rd_data_way1_out_56 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_57 <= 22'h0;
    end else if (_T_1512) begin
      btb_bank0_rd_data_way1_out_57 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_58 <= 22'h0;
    end else if (_T_1515) begin
      btb_bank0_rd_data_way1_out_58 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_59 <= 22'h0;
    end else if (_T_1518) begin
      btb_bank0_rd_data_way1_out_59 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_60 <= 22'h0;
    end else if (_T_1521) begin
      btb_bank0_rd_data_way1_out_60 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_61 <= 22'h0;
    end else if (_T_1524) begin
      btb_bank0_rd_data_way1_out_61 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_62 <= 22'h0;
    end else if (_T_1527) begin
      btb_bank0_rd_data_way1_out_62 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_63 <= 22'h0;
    end else if (_T_1530) begin
      btb_bank0_rd_data_way1_out_63 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_64 <= 22'h0;
    end else if (_T_1533) begin
      btb_bank0_rd_data_way1_out_64 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_65 <= 22'h0;
    end else if (_T_1536) begin
      btb_bank0_rd_data_way1_out_65 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_66 <= 22'h0;
    end else if (_T_1539) begin
      btb_bank0_rd_data_way1_out_66 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_67 <= 22'h0;
    end else if (_T_1542) begin
      btb_bank0_rd_data_way1_out_67 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_68 <= 22'h0;
    end else if (_T_1545) begin
      btb_bank0_rd_data_way1_out_68 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_69 <= 22'h0;
    end else if (_T_1548) begin
      btb_bank0_rd_data_way1_out_69 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_70 <= 22'h0;
    end else if (_T_1551) begin
      btb_bank0_rd_data_way1_out_70 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_71 <= 22'h0;
    end else if (_T_1554) begin
      btb_bank0_rd_data_way1_out_71 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_72 <= 22'h0;
    end else if (_T_1557) begin
      btb_bank0_rd_data_way1_out_72 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_73 <= 22'h0;
    end else if (_T_1560) begin
      btb_bank0_rd_data_way1_out_73 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_74 <= 22'h0;
    end else if (_T_1563) begin
      btb_bank0_rd_data_way1_out_74 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_75 <= 22'h0;
    end else if (_T_1566) begin
      btb_bank0_rd_data_way1_out_75 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_76 <= 22'h0;
    end else if (_T_1569) begin
      btb_bank0_rd_data_way1_out_76 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_77 <= 22'h0;
    end else if (_T_1572) begin
      btb_bank0_rd_data_way1_out_77 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_78 <= 22'h0;
    end else if (_T_1575) begin
      btb_bank0_rd_data_way1_out_78 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_79 <= 22'h0;
    end else if (_T_1578) begin
      btb_bank0_rd_data_way1_out_79 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_80 <= 22'h0;
    end else if (_T_1581) begin
      btb_bank0_rd_data_way1_out_80 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_81 <= 22'h0;
    end else if (_T_1584) begin
      btb_bank0_rd_data_way1_out_81 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_82 <= 22'h0;
    end else if (_T_1587) begin
      btb_bank0_rd_data_way1_out_82 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_83 <= 22'h0;
    end else if (_T_1590) begin
      btb_bank0_rd_data_way1_out_83 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_84 <= 22'h0;
    end else if (_T_1593) begin
      btb_bank0_rd_data_way1_out_84 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_85 <= 22'h0;
    end else if (_T_1596) begin
      btb_bank0_rd_data_way1_out_85 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_86 <= 22'h0;
    end else if (_T_1599) begin
      btb_bank0_rd_data_way1_out_86 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_87 <= 22'h0;
    end else if (_T_1602) begin
      btb_bank0_rd_data_way1_out_87 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_88 <= 22'h0;
    end else if (_T_1605) begin
      btb_bank0_rd_data_way1_out_88 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_89 <= 22'h0;
    end else if (_T_1608) begin
      btb_bank0_rd_data_way1_out_89 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_90 <= 22'h0;
    end else if (_T_1611) begin
      btb_bank0_rd_data_way1_out_90 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_91 <= 22'h0;
    end else if (_T_1614) begin
      btb_bank0_rd_data_way1_out_91 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_92 <= 22'h0;
    end else if (_T_1617) begin
      btb_bank0_rd_data_way1_out_92 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_93 <= 22'h0;
    end else if (_T_1620) begin
      btb_bank0_rd_data_way1_out_93 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_94 <= 22'h0;
    end else if (_T_1623) begin
      btb_bank0_rd_data_way1_out_94 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_95 <= 22'h0;
    end else if (_T_1626) begin
      btb_bank0_rd_data_way1_out_95 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_96 <= 22'h0;
    end else if (_T_1629) begin
      btb_bank0_rd_data_way1_out_96 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_97 <= 22'h0;
    end else if (_T_1632) begin
      btb_bank0_rd_data_way1_out_97 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_98 <= 22'h0;
    end else if (_T_1635) begin
      btb_bank0_rd_data_way1_out_98 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_99 <= 22'h0;
    end else if (_T_1638) begin
      btb_bank0_rd_data_way1_out_99 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_100 <= 22'h0;
    end else if (_T_1641) begin
      btb_bank0_rd_data_way1_out_100 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_101 <= 22'h0;
    end else if (_T_1644) begin
      btb_bank0_rd_data_way1_out_101 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_102 <= 22'h0;
    end else if (_T_1647) begin
      btb_bank0_rd_data_way1_out_102 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_103 <= 22'h0;
    end else if (_T_1650) begin
      btb_bank0_rd_data_way1_out_103 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_104 <= 22'h0;
    end else if (_T_1653) begin
      btb_bank0_rd_data_way1_out_104 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_105 <= 22'h0;
    end else if (_T_1656) begin
      btb_bank0_rd_data_way1_out_105 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_106 <= 22'h0;
    end else if (_T_1659) begin
      btb_bank0_rd_data_way1_out_106 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_107 <= 22'h0;
    end else if (_T_1662) begin
      btb_bank0_rd_data_way1_out_107 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_108 <= 22'h0;
    end else if (_T_1665) begin
      btb_bank0_rd_data_way1_out_108 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_109 <= 22'h0;
    end else if (_T_1668) begin
      btb_bank0_rd_data_way1_out_109 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_110 <= 22'h0;
    end else if (_T_1671) begin
      btb_bank0_rd_data_way1_out_110 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_111 <= 22'h0;
    end else if (_T_1674) begin
      btb_bank0_rd_data_way1_out_111 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_112 <= 22'h0;
    end else if (_T_1677) begin
      btb_bank0_rd_data_way1_out_112 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_113 <= 22'h0;
    end else if (_T_1680) begin
      btb_bank0_rd_data_way1_out_113 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_114 <= 22'h0;
    end else if (_T_1683) begin
      btb_bank0_rd_data_way1_out_114 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_115 <= 22'h0;
    end else if (_T_1686) begin
      btb_bank0_rd_data_way1_out_115 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_116 <= 22'h0;
    end else if (_T_1689) begin
      btb_bank0_rd_data_way1_out_116 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_117 <= 22'h0;
    end else if (_T_1692) begin
      btb_bank0_rd_data_way1_out_117 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_118 <= 22'h0;
    end else if (_T_1695) begin
      btb_bank0_rd_data_way1_out_118 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_119 <= 22'h0;
    end else if (_T_1698) begin
      btb_bank0_rd_data_way1_out_119 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_120 <= 22'h0;
    end else if (_T_1701) begin
      btb_bank0_rd_data_way1_out_120 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_121 <= 22'h0;
    end else if (_T_1704) begin
      btb_bank0_rd_data_way1_out_121 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_122 <= 22'h0;
    end else if (_T_1707) begin
      btb_bank0_rd_data_way1_out_122 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_123 <= 22'h0;
    end else if (_T_1710) begin
      btb_bank0_rd_data_way1_out_123 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_124 <= 22'h0;
    end else if (_T_1713) begin
      btb_bank0_rd_data_way1_out_124 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_125 <= 22'h0;
    end else if (_T_1716) begin
      btb_bank0_rd_data_way1_out_125 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_126 <= 22'h0;
    end else if (_T_1719) begin
      btb_bank0_rd_data_way1_out_126 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_127 <= 22'h0;
    end else if (_T_1722) begin
      btb_bank0_rd_data_way1_out_127 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_128 <= 22'h0;
    end else if (_T_1725) begin
      btb_bank0_rd_data_way1_out_128 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_129 <= 22'h0;
    end else if (_T_1728) begin
      btb_bank0_rd_data_way1_out_129 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_130 <= 22'h0;
    end else if (_T_1731) begin
      btb_bank0_rd_data_way1_out_130 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_131 <= 22'h0;
    end else if (_T_1734) begin
      btb_bank0_rd_data_way1_out_131 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_132 <= 22'h0;
    end else if (_T_1737) begin
      btb_bank0_rd_data_way1_out_132 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_133 <= 22'h0;
    end else if (_T_1740) begin
      btb_bank0_rd_data_way1_out_133 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_134 <= 22'h0;
    end else if (_T_1743) begin
      btb_bank0_rd_data_way1_out_134 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_135 <= 22'h0;
    end else if (_T_1746) begin
      btb_bank0_rd_data_way1_out_135 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_136 <= 22'h0;
    end else if (_T_1749) begin
      btb_bank0_rd_data_way1_out_136 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_137 <= 22'h0;
    end else if (_T_1752) begin
      btb_bank0_rd_data_way1_out_137 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_138 <= 22'h0;
    end else if (_T_1755) begin
      btb_bank0_rd_data_way1_out_138 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_139 <= 22'h0;
    end else if (_T_1758) begin
      btb_bank0_rd_data_way1_out_139 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_140 <= 22'h0;
    end else if (_T_1761) begin
      btb_bank0_rd_data_way1_out_140 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_141 <= 22'h0;
    end else if (_T_1764) begin
      btb_bank0_rd_data_way1_out_141 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_142 <= 22'h0;
    end else if (_T_1767) begin
      btb_bank0_rd_data_way1_out_142 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_143 <= 22'h0;
    end else if (_T_1770) begin
      btb_bank0_rd_data_way1_out_143 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_144 <= 22'h0;
    end else if (_T_1773) begin
      btb_bank0_rd_data_way1_out_144 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_145 <= 22'h0;
    end else if (_T_1776) begin
      btb_bank0_rd_data_way1_out_145 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_146 <= 22'h0;
    end else if (_T_1779) begin
      btb_bank0_rd_data_way1_out_146 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_147 <= 22'h0;
    end else if (_T_1782) begin
      btb_bank0_rd_data_way1_out_147 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_148 <= 22'h0;
    end else if (_T_1785) begin
      btb_bank0_rd_data_way1_out_148 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_149 <= 22'h0;
    end else if (_T_1788) begin
      btb_bank0_rd_data_way1_out_149 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_150 <= 22'h0;
    end else if (_T_1791) begin
      btb_bank0_rd_data_way1_out_150 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_151 <= 22'h0;
    end else if (_T_1794) begin
      btb_bank0_rd_data_way1_out_151 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_152 <= 22'h0;
    end else if (_T_1797) begin
      btb_bank0_rd_data_way1_out_152 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_153 <= 22'h0;
    end else if (_T_1800) begin
      btb_bank0_rd_data_way1_out_153 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_154 <= 22'h0;
    end else if (_T_1803) begin
      btb_bank0_rd_data_way1_out_154 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_155 <= 22'h0;
    end else if (_T_1806) begin
      btb_bank0_rd_data_way1_out_155 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_156 <= 22'h0;
    end else if (_T_1809) begin
      btb_bank0_rd_data_way1_out_156 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_157 <= 22'h0;
    end else if (_T_1812) begin
      btb_bank0_rd_data_way1_out_157 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_158 <= 22'h0;
    end else if (_T_1815) begin
      btb_bank0_rd_data_way1_out_158 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_159 <= 22'h0;
    end else if (_T_1818) begin
      btb_bank0_rd_data_way1_out_159 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_160 <= 22'h0;
    end else if (_T_1821) begin
      btb_bank0_rd_data_way1_out_160 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_161 <= 22'h0;
    end else if (_T_1824) begin
      btb_bank0_rd_data_way1_out_161 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_162 <= 22'h0;
    end else if (_T_1827) begin
      btb_bank0_rd_data_way1_out_162 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_163 <= 22'h0;
    end else if (_T_1830) begin
      btb_bank0_rd_data_way1_out_163 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_164 <= 22'h0;
    end else if (_T_1833) begin
      btb_bank0_rd_data_way1_out_164 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_165 <= 22'h0;
    end else if (_T_1836) begin
      btb_bank0_rd_data_way1_out_165 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_166 <= 22'h0;
    end else if (_T_1839) begin
      btb_bank0_rd_data_way1_out_166 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_167 <= 22'h0;
    end else if (_T_1842) begin
      btb_bank0_rd_data_way1_out_167 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_168 <= 22'h0;
    end else if (_T_1845) begin
      btb_bank0_rd_data_way1_out_168 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_169 <= 22'h0;
    end else if (_T_1848) begin
      btb_bank0_rd_data_way1_out_169 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_170 <= 22'h0;
    end else if (_T_1851) begin
      btb_bank0_rd_data_way1_out_170 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_171 <= 22'h0;
    end else if (_T_1854) begin
      btb_bank0_rd_data_way1_out_171 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_172 <= 22'h0;
    end else if (_T_1857) begin
      btb_bank0_rd_data_way1_out_172 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_173 <= 22'h0;
    end else if (_T_1860) begin
      btb_bank0_rd_data_way1_out_173 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_174 <= 22'h0;
    end else if (_T_1863) begin
      btb_bank0_rd_data_way1_out_174 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_175 <= 22'h0;
    end else if (_T_1866) begin
      btb_bank0_rd_data_way1_out_175 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_176 <= 22'h0;
    end else if (_T_1869) begin
      btb_bank0_rd_data_way1_out_176 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_177 <= 22'h0;
    end else if (_T_1872) begin
      btb_bank0_rd_data_way1_out_177 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_178 <= 22'h0;
    end else if (_T_1875) begin
      btb_bank0_rd_data_way1_out_178 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_179 <= 22'h0;
    end else if (_T_1878) begin
      btb_bank0_rd_data_way1_out_179 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_180 <= 22'h0;
    end else if (_T_1881) begin
      btb_bank0_rd_data_way1_out_180 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_181 <= 22'h0;
    end else if (_T_1884) begin
      btb_bank0_rd_data_way1_out_181 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_182 <= 22'h0;
    end else if (_T_1887) begin
      btb_bank0_rd_data_way1_out_182 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_183 <= 22'h0;
    end else if (_T_1890) begin
      btb_bank0_rd_data_way1_out_183 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_184 <= 22'h0;
    end else if (_T_1893) begin
      btb_bank0_rd_data_way1_out_184 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_185 <= 22'h0;
    end else if (_T_1896) begin
      btb_bank0_rd_data_way1_out_185 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_186 <= 22'h0;
    end else if (_T_1899) begin
      btb_bank0_rd_data_way1_out_186 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_187 <= 22'h0;
    end else if (_T_1902) begin
      btb_bank0_rd_data_way1_out_187 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_188 <= 22'h0;
    end else if (_T_1905) begin
      btb_bank0_rd_data_way1_out_188 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_189 <= 22'h0;
    end else if (_T_1908) begin
      btb_bank0_rd_data_way1_out_189 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_190 <= 22'h0;
    end else if (_T_1911) begin
      btb_bank0_rd_data_way1_out_190 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_191 <= 22'h0;
    end else if (_T_1914) begin
      btb_bank0_rd_data_way1_out_191 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_192 <= 22'h0;
    end else if (_T_1917) begin
      btb_bank0_rd_data_way1_out_192 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_193 <= 22'h0;
    end else if (_T_1920) begin
      btb_bank0_rd_data_way1_out_193 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_194 <= 22'h0;
    end else if (_T_1923) begin
      btb_bank0_rd_data_way1_out_194 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_195 <= 22'h0;
    end else if (_T_1926) begin
      btb_bank0_rd_data_way1_out_195 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_196 <= 22'h0;
    end else if (_T_1929) begin
      btb_bank0_rd_data_way1_out_196 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_197 <= 22'h0;
    end else if (_T_1932) begin
      btb_bank0_rd_data_way1_out_197 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_198 <= 22'h0;
    end else if (_T_1935) begin
      btb_bank0_rd_data_way1_out_198 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_199 <= 22'h0;
    end else if (_T_1938) begin
      btb_bank0_rd_data_way1_out_199 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_200 <= 22'h0;
    end else if (_T_1941) begin
      btb_bank0_rd_data_way1_out_200 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_201 <= 22'h0;
    end else if (_T_1944) begin
      btb_bank0_rd_data_way1_out_201 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_202 <= 22'h0;
    end else if (_T_1947) begin
      btb_bank0_rd_data_way1_out_202 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_203 <= 22'h0;
    end else if (_T_1950) begin
      btb_bank0_rd_data_way1_out_203 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_204 <= 22'h0;
    end else if (_T_1953) begin
      btb_bank0_rd_data_way1_out_204 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_205 <= 22'h0;
    end else if (_T_1956) begin
      btb_bank0_rd_data_way1_out_205 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_206 <= 22'h0;
    end else if (_T_1959) begin
      btb_bank0_rd_data_way1_out_206 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_207 <= 22'h0;
    end else if (_T_1962) begin
      btb_bank0_rd_data_way1_out_207 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_208 <= 22'h0;
    end else if (_T_1965) begin
      btb_bank0_rd_data_way1_out_208 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_209 <= 22'h0;
    end else if (_T_1968) begin
      btb_bank0_rd_data_way1_out_209 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_210 <= 22'h0;
    end else if (_T_1971) begin
      btb_bank0_rd_data_way1_out_210 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_211 <= 22'h0;
    end else if (_T_1974) begin
      btb_bank0_rd_data_way1_out_211 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_212 <= 22'h0;
    end else if (_T_1977) begin
      btb_bank0_rd_data_way1_out_212 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_213 <= 22'h0;
    end else if (_T_1980) begin
      btb_bank0_rd_data_way1_out_213 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_214 <= 22'h0;
    end else if (_T_1983) begin
      btb_bank0_rd_data_way1_out_214 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_215 <= 22'h0;
    end else if (_T_1986) begin
      btb_bank0_rd_data_way1_out_215 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_216 <= 22'h0;
    end else if (_T_1989) begin
      btb_bank0_rd_data_way1_out_216 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_217 <= 22'h0;
    end else if (_T_1992) begin
      btb_bank0_rd_data_way1_out_217 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_218 <= 22'h0;
    end else if (_T_1995) begin
      btb_bank0_rd_data_way1_out_218 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_219 <= 22'h0;
    end else if (_T_1998) begin
      btb_bank0_rd_data_way1_out_219 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_220 <= 22'h0;
    end else if (_T_2001) begin
      btb_bank0_rd_data_way1_out_220 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_221 <= 22'h0;
    end else if (_T_2004) begin
      btb_bank0_rd_data_way1_out_221 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_222 <= 22'h0;
    end else if (_T_2007) begin
      btb_bank0_rd_data_way1_out_222 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_223 <= 22'h0;
    end else if (_T_2010) begin
      btb_bank0_rd_data_way1_out_223 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_224 <= 22'h0;
    end else if (_T_2013) begin
      btb_bank0_rd_data_way1_out_224 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_225 <= 22'h0;
    end else if (_T_2016) begin
      btb_bank0_rd_data_way1_out_225 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_226 <= 22'h0;
    end else if (_T_2019) begin
      btb_bank0_rd_data_way1_out_226 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_227 <= 22'h0;
    end else if (_T_2022) begin
      btb_bank0_rd_data_way1_out_227 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_228 <= 22'h0;
    end else if (_T_2025) begin
      btb_bank0_rd_data_way1_out_228 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_229 <= 22'h0;
    end else if (_T_2028) begin
      btb_bank0_rd_data_way1_out_229 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_230 <= 22'h0;
    end else if (_T_2031) begin
      btb_bank0_rd_data_way1_out_230 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_231 <= 22'h0;
    end else if (_T_2034) begin
      btb_bank0_rd_data_way1_out_231 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_232 <= 22'h0;
    end else if (_T_2037) begin
      btb_bank0_rd_data_way1_out_232 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_233 <= 22'h0;
    end else if (_T_2040) begin
      btb_bank0_rd_data_way1_out_233 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_234 <= 22'h0;
    end else if (_T_2043) begin
      btb_bank0_rd_data_way1_out_234 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_235 <= 22'h0;
    end else if (_T_2046) begin
      btb_bank0_rd_data_way1_out_235 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_236 <= 22'h0;
    end else if (_T_2049) begin
      btb_bank0_rd_data_way1_out_236 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_237 <= 22'h0;
    end else if (_T_2052) begin
      btb_bank0_rd_data_way1_out_237 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_238 <= 22'h0;
    end else if (_T_2055) begin
      btb_bank0_rd_data_way1_out_238 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_239 <= 22'h0;
    end else if (_T_2058) begin
      btb_bank0_rd_data_way1_out_239 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_240 <= 22'h0;
    end else if (_T_2061) begin
      btb_bank0_rd_data_way1_out_240 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_241 <= 22'h0;
    end else if (_T_2064) begin
      btb_bank0_rd_data_way1_out_241 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_242 <= 22'h0;
    end else if (_T_2067) begin
      btb_bank0_rd_data_way1_out_242 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_243 <= 22'h0;
    end else if (_T_2070) begin
      btb_bank0_rd_data_way1_out_243 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_244 <= 22'h0;
    end else if (_T_2073) begin
      btb_bank0_rd_data_way1_out_244 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_245 <= 22'h0;
    end else if (_T_2076) begin
      btb_bank0_rd_data_way1_out_245 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_246 <= 22'h0;
    end else if (_T_2079) begin
      btb_bank0_rd_data_way1_out_246 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_247 <= 22'h0;
    end else if (_T_2082) begin
      btb_bank0_rd_data_way1_out_247 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_248 <= 22'h0;
    end else if (_T_2085) begin
      btb_bank0_rd_data_way1_out_248 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_249 <= 22'h0;
    end else if (_T_2088) begin
      btb_bank0_rd_data_way1_out_249 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_250 <= 22'h0;
    end else if (_T_2091) begin
      btb_bank0_rd_data_way1_out_250 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_251 <= 22'h0;
    end else if (_T_2094) begin
      btb_bank0_rd_data_way1_out_251 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_252 <= 22'h0;
    end else if (_T_2097) begin
      btb_bank0_rd_data_way1_out_252 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_253 <= 22'h0;
    end else if (_T_2100) begin
      btb_bank0_rd_data_way1_out_253 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_254 <= 22'h0;
    end else if (_T_2103) begin
      btb_bank0_rd_data_way1_out_254 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_255 <= 22'h0;
    end else if (_T_2106) begin
      btb_bank0_rd_data_way1_out_255 <= btb_wr_data;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fghr <= 8'h0;
    end else begin
      fghr <= _T_337 | _T_336;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_0 <= 2'h0;
    end else if (bht_bank_sel_1_0_0) begin
      if (_T_8802) begin
        bht_bank_rd_data_out_1_0 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_0 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_1 <= 2'h0;
    end else if (bht_bank_sel_1_0_1) begin
      if (_T_8811) begin
        bht_bank_rd_data_out_1_1 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_1 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_2 <= 2'h0;
    end else if (bht_bank_sel_1_0_2) begin
      if (_T_8820) begin
        bht_bank_rd_data_out_1_2 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_2 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_3 <= 2'h0;
    end else if (bht_bank_sel_1_0_3) begin
      if (_T_8829) begin
        bht_bank_rd_data_out_1_3 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_3 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_4 <= 2'h0;
    end else if (bht_bank_sel_1_0_4) begin
      if (_T_8838) begin
        bht_bank_rd_data_out_1_4 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_4 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_5 <= 2'h0;
    end else if (bht_bank_sel_1_0_5) begin
      if (_T_8847) begin
        bht_bank_rd_data_out_1_5 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_5 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_6 <= 2'h0;
    end else if (bht_bank_sel_1_0_6) begin
      if (_T_8856) begin
        bht_bank_rd_data_out_1_6 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_6 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_7 <= 2'h0;
    end else if (bht_bank_sel_1_0_7) begin
      if (_T_8865) begin
        bht_bank_rd_data_out_1_7 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_7 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_8 <= 2'h0;
    end else if (bht_bank_sel_1_0_8) begin
      if (_T_8874) begin
        bht_bank_rd_data_out_1_8 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_8 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_9 <= 2'h0;
    end else if (bht_bank_sel_1_0_9) begin
      if (_T_8883) begin
        bht_bank_rd_data_out_1_9 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_9 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_10 <= 2'h0;
    end else if (bht_bank_sel_1_0_10) begin
      if (_T_8892) begin
        bht_bank_rd_data_out_1_10 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_10 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_11 <= 2'h0;
    end else if (bht_bank_sel_1_0_11) begin
      if (_T_8901) begin
        bht_bank_rd_data_out_1_11 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_11 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_12 <= 2'h0;
    end else if (bht_bank_sel_1_0_12) begin
      if (_T_8910) begin
        bht_bank_rd_data_out_1_12 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_12 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_13 <= 2'h0;
    end else if (bht_bank_sel_1_0_13) begin
      if (_T_8919) begin
        bht_bank_rd_data_out_1_13 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_13 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_14 <= 2'h0;
    end else if (bht_bank_sel_1_0_14) begin
      if (_T_8928) begin
        bht_bank_rd_data_out_1_14 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_14 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_15 <= 2'h0;
    end else if (bht_bank_sel_1_0_15) begin
      if (_T_8937) begin
        bht_bank_rd_data_out_1_15 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_15 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_16 <= 2'h0;
    end else if (bht_bank_sel_1_1_0) begin
      if (_T_8946) begin
        bht_bank_rd_data_out_1_16 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_16 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_17 <= 2'h0;
    end else if (bht_bank_sel_1_1_1) begin
      if (_T_8955) begin
        bht_bank_rd_data_out_1_17 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_17 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_18 <= 2'h0;
    end else if (bht_bank_sel_1_1_2) begin
      if (_T_8964) begin
        bht_bank_rd_data_out_1_18 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_18 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_19 <= 2'h0;
    end else if (bht_bank_sel_1_1_3) begin
      if (_T_8973) begin
        bht_bank_rd_data_out_1_19 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_19 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_20 <= 2'h0;
    end else if (bht_bank_sel_1_1_4) begin
      if (_T_8982) begin
        bht_bank_rd_data_out_1_20 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_20 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_21 <= 2'h0;
    end else if (bht_bank_sel_1_1_5) begin
      if (_T_8991) begin
        bht_bank_rd_data_out_1_21 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_21 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_22 <= 2'h0;
    end else if (bht_bank_sel_1_1_6) begin
      if (_T_9000) begin
        bht_bank_rd_data_out_1_22 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_22 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_23 <= 2'h0;
    end else if (bht_bank_sel_1_1_7) begin
      if (_T_9009) begin
        bht_bank_rd_data_out_1_23 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_23 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_24 <= 2'h0;
    end else if (bht_bank_sel_1_1_8) begin
      if (_T_9018) begin
        bht_bank_rd_data_out_1_24 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_24 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_25 <= 2'h0;
    end else if (bht_bank_sel_1_1_9) begin
      if (_T_9027) begin
        bht_bank_rd_data_out_1_25 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_25 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_26 <= 2'h0;
    end else if (bht_bank_sel_1_1_10) begin
      if (_T_9036) begin
        bht_bank_rd_data_out_1_26 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_26 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_27 <= 2'h0;
    end else if (bht_bank_sel_1_1_11) begin
      if (_T_9045) begin
        bht_bank_rd_data_out_1_27 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_27 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_28 <= 2'h0;
    end else if (bht_bank_sel_1_1_12) begin
      if (_T_9054) begin
        bht_bank_rd_data_out_1_28 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_28 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_29 <= 2'h0;
    end else if (bht_bank_sel_1_1_13) begin
      if (_T_9063) begin
        bht_bank_rd_data_out_1_29 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_29 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_30 <= 2'h0;
    end else if (bht_bank_sel_1_1_14) begin
      if (_T_9072) begin
        bht_bank_rd_data_out_1_30 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_30 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_31 <= 2'h0;
    end else if (bht_bank_sel_1_1_15) begin
      if (_T_9081) begin
        bht_bank_rd_data_out_1_31 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_31 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_32 <= 2'h0;
    end else if (bht_bank_sel_1_2_0) begin
      if (_T_9090) begin
        bht_bank_rd_data_out_1_32 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_32 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_33 <= 2'h0;
    end else if (bht_bank_sel_1_2_1) begin
      if (_T_9099) begin
        bht_bank_rd_data_out_1_33 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_33 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_34 <= 2'h0;
    end else if (bht_bank_sel_1_2_2) begin
      if (_T_9108) begin
        bht_bank_rd_data_out_1_34 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_34 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_35 <= 2'h0;
    end else if (bht_bank_sel_1_2_3) begin
      if (_T_9117) begin
        bht_bank_rd_data_out_1_35 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_35 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_36 <= 2'h0;
    end else if (bht_bank_sel_1_2_4) begin
      if (_T_9126) begin
        bht_bank_rd_data_out_1_36 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_36 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_37 <= 2'h0;
    end else if (bht_bank_sel_1_2_5) begin
      if (_T_9135) begin
        bht_bank_rd_data_out_1_37 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_37 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_38 <= 2'h0;
    end else if (bht_bank_sel_1_2_6) begin
      if (_T_9144) begin
        bht_bank_rd_data_out_1_38 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_38 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_39 <= 2'h0;
    end else if (bht_bank_sel_1_2_7) begin
      if (_T_9153) begin
        bht_bank_rd_data_out_1_39 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_39 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_40 <= 2'h0;
    end else if (bht_bank_sel_1_2_8) begin
      if (_T_9162) begin
        bht_bank_rd_data_out_1_40 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_40 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_41 <= 2'h0;
    end else if (bht_bank_sel_1_2_9) begin
      if (_T_9171) begin
        bht_bank_rd_data_out_1_41 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_41 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_42 <= 2'h0;
    end else if (bht_bank_sel_1_2_10) begin
      if (_T_9180) begin
        bht_bank_rd_data_out_1_42 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_42 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_43 <= 2'h0;
    end else if (bht_bank_sel_1_2_11) begin
      if (_T_9189) begin
        bht_bank_rd_data_out_1_43 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_43 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_44 <= 2'h0;
    end else if (bht_bank_sel_1_2_12) begin
      if (_T_9198) begin
        bht_bank_rd_data_out_1_44 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_44 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_45 <= 2'h0;
    end else if (bht_bank_sel_1_2_13) begin
      if (_T_9207) begin
        bht_bank_rd_data_out_1_45 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_45 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_46 <= 2'h0;
    end else if (bht_bank_sel_1_2_14) begin
      if (_T_9216) begin
        bht_bank_rd_data_out_1_46 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_46 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_47 <= 2'h0;
    end else if (bht_bank_sel_1_2_15) begin
      if (_T_9225) begin
        bht_bank_rd_data_out_1_47 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_47 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_48 <= 2'h0;
    end else if (bht_bank_sel_1_3_0) begin
      if (_T_9234) begin
        bht_bank_rd_data_out_1_48 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_48 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_49 <= 2'h0;
    end else if (bht_bank_sel_1_3_1) begin
      if (_T_9243) begin
        bht_bank_rd_data_out_1_49 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_49 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_50 <= 2'h0;
    end else if (bht_bank_sel_1_3_2) begin
      if (_T_9252) begin
        bht_bank_rd_data_out_1_50 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_50 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_51 <= 2'h0;
    end else if (bht_bank_sel_1_3_3) begin
      if (_T_9261) begin
        bht_bank_rd_data_out_1_51 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_51 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_52 <= 2'h0;
    end else if (bht_bank_sel_1_3_4) begin
      if (_T_9270) begin
        bht_bank_rd_data_out_1_52 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_52 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_53 <= 2'h0;
    end else if (bht_bank_sel_1_3_5) begin
      if (_T_9279) begin
        bht_bank_rd_data_out_1_53 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_53 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_54 <= 2'h0;
    end else if (bht_bank_sel_1_3_6) begin
      if (_T_9288) begin
        bht_bank_rd_data_out_1_54 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_54 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_55 <= 2'h0;
    end else if (bht_bank_sel_1_3_7) begin
      if (_T_9297) begin
        bht_bank_rd_data_out_1_55 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_55 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_56 <= 2'h0;
    end else if (bht_bank_sel_1_3_8) begin
      if (_T_9306) begin
        bht_bank_rd_data_out_1_56 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_56 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_57 <= 2'h0;
    end else if (bht_bank_sel_1_3_9) begin
      if (_T_9315) begin
        bht_bank_rd_data_out_1_57 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_57 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_58 <= 2'h0;
    end else if (bht_bank_sel_1_3_10) begin
      if (_T_9324) begin
        bht_bank_rd_data_out_1_58 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_58 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_59 <= 2'h0;
    end else if (bht_bank_sel_1_3_11) begin
      if (_T_9333) begin
        bht_bank_rd_data_out_1_59 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_59 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_60 <= 2'h0;
    end else if (bht_bank_sel_1_3_12) begin
      if (_T_9342) begin
        bht_bank_rd_data_out_1_60 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_60 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_61 <= 2'h0;
    end else if (bht_bank_sel_1_3_13) begin
      if (_T_9351) begin
        bht_bank_rd_data_out_1_61 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_61 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_62 <= 2'h0;
    end else if (bht_bank_sel_1_3_14) begin
      if (_T_9360) begin
        bht_bank_rd_data_out_1_62 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_62 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_63 <= 2'h0;
    end else if (bht_bank_sel_1_3_15) begin
      if (_T_9369) begin
        bht_bank_rd_data_out_1_63 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_63 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_64 <= 2'h0;
    end else if (bht_bank_sel_1_4_0) begin
      if (_T_9378) begin
        bht_bank_rd_data_out_1_64 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_64 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_65 <= 2'h0;
    end else if (bht_bank_sel_1_4_1) begin
      if (_T_9387) begin
        bht_bank_rd_data_out_1_65 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_65 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_66 <= 2'h0;
    end else if (bht_bank_sel_1_4_2) begin
      if (_T_9396) begin
        bht_bank_rd_data_out_1_66 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_66 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_67 <= 2'h0;
    end else if (bht_bank_sel_1_4_3) begin
      if (_T_9405) begin
        bht_bank_rd_data_out_1_67 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_67 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_68 <= 2'h0;
    end else if (bht_bank_sel_1_4_4) begin
      if (_T_9414) begin
        bht_bank_rd_data_out_1_68 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_68 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_69 <= 2'h0;
    end else if (bht_bank_sel_1_4_5) begin
      if (_T_9423) begin
        bht_bank_rd_data_out_1_69 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_69 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_70 <= 2'h0;
    end else if (bht_bank_sel_1_4_6) begin
      if (_T_9432) begin
        bht_bank_rd_data_out_1_70 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_70 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_71 <= 2'h0;
    end else if (bht_bank_sel_1_4_7) begin
      if (_T_9441) begin
        bht_bank_rd_data_out_1_71 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_71 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_72 <= 2'h0;
    end else if (bht_bank_sel_1_4_8) begin
      if (_T_9450) begin
        bht_bank_rd_data_out_1_72 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_72 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_73 <= 2'h0;
    end else if (bht_bank_sel_1_4_9) begin
      if (_T_9459) begin
        bht_bank_rd_data_out_1_73 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_73 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_74 <= 2'h0;
    end else if (bht_bank_sel_1_4_10) begin
      if (_T_9468) begin
        bht_bank_rd_data_out_1_74 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_74 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_75 <= 2'h0;
    end else if (bht_bank_sel_1_4_11) begin
      if (_T_9477) begin
        bht_bank_rd_data_out_1_75 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_75 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_76 <= 2'h0;
    end else if (bht_bank_sel_1_4_12) begin
      if (_T_9486) begin
        bht_bank_rd_data_out_1_76 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_76 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_77 <= 2'h0;
    end else if (bht_bank_sel_1_4_13) begin
      if (_T_9495) begin
        bht_bank_rd_data_out_1_77 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_77 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_78 <= 2'h0;
    end else if (bht_bank_sel_1_4_14) begin
      if (_T_9504) begin
        bht_bank_rd_data_out_1_78 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_78 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_79 <= 2'h0;
    end else if (bht_bank_sel_1_4_15) begin
      if (_T_9513) begin
        bht_bank_rd_data_out_1_79 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_79 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_80 <= 2'h0;
    end else if (bht_bank_sel_1_5_0) begin
      if (_T_9522) begin
        bht_bank_rd_data_out_1_80 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_80 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_81 <= 2'h0;
    end else if (bht_bank_sel_1_5_1) begin
      if (_T_9531) begin
        bht_bank_rd_data_out_1_81 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_81 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_82 <= 2'h0;
    end else if (bht_bank_sel_1_5_2) begin
      if (_T_9540) begin
        bht_bank_rd_data_out_1_82 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_82 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_83 <= 2'h0;
    end else if (bht_bank_sel_1_5_3) begin
      if (_T_9549) begin
        bht_bank_rd_data_out_1_83 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_83 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_84 <= 2'h0;
    end else if (bht_bank_sel_1_5_4) begin
      if (_T_9558) begin
        bht_bank_rd_data_out_1_84 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_84 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_85 <= 2'h0;
    end else if (bht_bank_sel_1_5_5) begin
      if (_T_9567) begin
        bht_bank_rd_data_out_1_85 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_85 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_86 <= 2'h0;
    end else if (bht_bank_sel_1_5_6) begin
      if (_T_9576) begin
        bht_bank_rd_data_out_1_86 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_86 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_87 <= 2'h0;
    end else if (bht_bank_sel_1_5_7) begin
      if (_T_9585) begin
        bht_bank_rd_data_out_1_87 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_87 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_88 <= 2'h0;
    end else if (bht_bank_sel_1_5_8) begin
      if (_T_9594) begin
        bht_bank_rd_data_out_1_88 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_88 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_89 <= 2'h0;
    end else if (bht_bank_sel_1_5_9) begin
      if (_T_9603) begin
        bht_bank_rd_data_out_1_89 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_89 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_90 <= 2'h0;
    end else if (bht_bank_sel_1_5_10) begin
      if (_T_9612) begin
        bht_bank_rd_data_out_1_90 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_90 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_91 <= 2'h0;
    end else if (bht_bank_sel_1_5_11) begin
      if (_T_9621) begin
        bht_bank_rd_data_out_1_91 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_91 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_92 <= 2'h0;
    end else if (bht_bank_sel_1_5_12) begin
      if (_T_9630) begin
        bht_bank_rd_data_out_1_92 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_92 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_93 <= 2'h0;
    end else if (bht_bank_sel_1_5_13) begin
      if (_T_9639) begin
        bht_bank_rd_data_out_1_93 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_93 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_94 <= 2'h0;
    end else if (bht_bank_sel_1_5_14) begin
      if (_T_9648) begin
        bht_bank_rd_data_out_1_94 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_94 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_95 <= 2'h0;
    end else if (bht_bank_sel_1_5_15) begin
      if (_T_9657) begin
        bht_bank_rd_data_out_1_95 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_95 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_96 <= 2'h0;
    end else if (bht_bank_sel_1_6_0) begin
      if (_T_9666) begin
        bht_bank_rd_data_out_1_96 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_96 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_97 <= 2'h0;
    end else if (bht_bank_sel_1_6_1) begin
      if (_T_9675) begin
        bht_bank_rd_data_out_1_97 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_97 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_98 <= 2'h0;
    end else if (bht_bank_sel_1_6_2) begin
      if (_T_9684) begin
        bht_bank_rd_data_out_1_98 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_98 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_99 <= 2'h0;
    end else if (bht_bank_sel_1_6_3) begin
      if (_T_9693) begin
        bht_bank_rd_data_out_1_99 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_99 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_100 <= 2'h0;
    end else if (bht_bank_sel_1_6_4) begin
      if (_T_9702) begin
        bht_bank_rd_data_out_1_100 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_100 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_101 <= 2'h0;
    end else if (bht_bank_sel_1_6_5) begin
      if (_T_9711) begin
        bht_bank_rd_data_out_1_101 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_101 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_102 <= 2'h0;
    end else if (bht_bank_sel_1_6_6) begin
      if (_T_9720) begin
        bht_bank_rd_data_out_1_102 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_102 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_103 <= 2'h0;
    end else if (bht_bank_sel_1_6_7) begin
      if (_T_9729) begin
        bht_bank_rd_data_out_1_103 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_103 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_104 <= 2'h0;
    end else if (bht_bank_sel_1_6_8) begin
      if (_T_9738) begin
        bht_bank_rd_data_out_1_104 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_104 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_105 <= 2'h0;
    end else if (bht_bank_sel_1_6_9) begin
      if (_T_9747) begin
        bht_bank_rd_data_out_1_105 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_105 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_106 <= 2'h0;
    end else if (bht_bank_sel_1_6_10) begin
      if (_T_9756) begin
        bht_bank_rd_data_out_1_106 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_106 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_107 <= 2'h0;
    end else if (bht_bank_sel_1_6_11) begin
      if (_T_9765) begin
        bht_bank_rd_data_out_1_107 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_107 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_108 <= 2'h0;
    end else if (bht_bank_sel_1_6_12) begin
      if (_T_9774) begin
        bht_bank_rd_data_out_1_108 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_108 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_109 <= 2'h0;
    end else if (bht_bank_sel_1_6_13) begin
      if (_T_9783) begin
        bht_bank_rd_data_out_1_109 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_109 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_110 <= 2'h0;
    end else if (bht_bank_sel_1_6_14) begin
      if (_T_9792) begin
        bht_bank_rd_data_out_1_110 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_110 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_111 <= 2'h0;
    end else if (bht_bank_sel_1_6_15) begin
      if (_T_9801) begin
        bht_bank_rd_data_out_1_111 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_111 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_112 <= 2'h0;
    end else if (bht_bank_sel_1_7_0) begin
      if (_T_9810) begin
        bht_bank_rd_data_out_1_112 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_112 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_113 <= 2'h0;
    end else if (bht_bank_sel_1_7_1) begin
      if (_T_9819) begin
        bht_bank_rd_data_out_1_113 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_113 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_114 <= 2'h0;
    end else if (bht_bank_sel_1_7_2) begin
      if (_T_9828) begin
        bht_bank_rd_data_out_1_114 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_114 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_115 <= 2'h0;
    end else if (bht_bank_sel_1_7_3) begin
      if (_T_9837) begin
        bht_bank_rd_data_out_1_115 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_115 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_116 <= 2'h0;
    end else if (bht_bank_sel_1_7_4) begin
      if (_T_9846) begin
        bht_bank_rd_data_out_1_116 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_116 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_117 <= 2'h0;
    end else if (bht_bank_sel_1_7_5) begin
      if (_T_9855) begin
        bht_bank_rd_data_out_1_117 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_117 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_118 <= 2'h0;
    end else if (bht_bank_sel_1_7_6) begin
      if (_T_9864) begin
        bht_bank_rd_data_out_1_118 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_118 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_119 <= 2'h0;
    end else if (bht_bank_sel_1_7_7) begin
      if (_T_9873) begin
        bht_bank_rd_data_out_1_119 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_119 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_120 <= 2'h0;
    end else if (bht_bank_sel_1_7_8) begin
      if (_T_9882) begin
        bht_bank_rd_data_out_1_120 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_120 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_121 <= 2'h0;
    end else if (bht_bank_sel_1_7_9) begin
      if (_T_9891) begin
        bht_bank_rd_data_out_1_121 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_121 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_122 <= 2'h0;
    end else if (bht_bank_sel_1_7_10) begin
      if (_T_9900) begin
        bht_bank_rd_data_out_1_122 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_122 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_123 <= 2'h0;
    end else if (bht_bank_sel_1_7_11) begin
      if (_T_9909) begin
        bht_bank_rd_data_out_1_123 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_123 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_124 <= 2'h0;
    end else if (bht_bank_sel_1_7_12) begin
      if (_T_9918) begin
        bht_bank_rd_data_out_1_124 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_124 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_125 <= 2'h0;
    end else if (bht_bank_sel_1_7_13) begin
      if (_T_9927) begin
        bht_bank_rd_data_out_1_125 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_125 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_126 <= 2'h0;
    end else if (bht_bank_sel_1_7_14) begin
      if (_T_9936) begin
        bht_bank_rd_data_out_1_126 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_126 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_127 <= 2'h0;
    end else if (bht_bank_sel_1_7_15) begin
      if (_T_9945) begin
        bht_bank_rd_data_out_1_127 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_127 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_128 <= 2'h0;
    end else if (bht_bank_sel_1_8_0) begin
      if (_T_9954) begin
        bht_bank_rd_data_out_1_128 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_128 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_129 <= 2'h0;
    end else if (bht_bank_sel_1_8_1) begin
      if (_T_9963) begin
        bht_bank_rd_data_out_1_129 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_129 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_130 <= 2'h0;
    end else if (bht_bank_sel_1_8_2) begin
      if (_T_9972) begin
        bht_bank_rd_data_out_1_130 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_130 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_131 <= 2'h0;
    end else if (bht_bank_sel_1_8_3) begin
      if (_T_9981) begin
        bht_bank_rd_data_out_1_131 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_131 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_132 <= 2'h0;
    end else if (bht_bank_sel_1_8_4) begin
      if (_T_9990) begin
        bht_bank_rd_data_out_1_132 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_132 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_133 <= 2'h0;
    end else if (bht_bank_sel_1_8_5) begin
      if (_T_9999) begin
        bht_bank_rd_data_out_1_133 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_133 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_134 <= 2'h0;
    end else if (bht_bank_sel_1_8_6) begin
      if (_T_10008) begin
        bht_bank_rd_data_out_1_134 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_134 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_135 <= 2'h0;
    end else if (bht_bank_sel_1_8_7) begin
      if (_T_10017) begin
        bht_bank_rd_data_out_1_135 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_135 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_136 <= 2'h0;
    end else if (bht_bank_sel_1_8_8) begin
      if (_T_10026) begin
        bht_bank_rd_data_out_1_136 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_136 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_137 <= 2'h0;
    end else if (bht_bank_sel_1_8_9) begin
      if (_T_10035) begin
        bht_bank_rd_data_out_1_137 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_137 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_138 <= 2'h0;
    end else if (bht_bank_sel_1_8_10) begin
      if (_T_10044) begin
        bht_bank_rd_data_out_1_138 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_138 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_139 <= 2'h0;
    end else if (bht_bank_sel_1_8_11) begin
      if (_T_10053) begin
        bht_bank_rd_data_out_1_139 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_139 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_140 <= 2'h0;
    end else if (bht_bank_sel_1_8_12) begin
      if (_T_10062) begin
        bht_bank_rd_data_out_1_140 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_140 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_141 <= 2'h0;
    end else if (bht_bank_sel_1_8_13) begin
      if (_T_10071) begin
        bht_bank_rd_data_out_1_141 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_141 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_142 <= 2'h0;
    end else if (bht_bank_sel_1_8_14) begin
      if (_T_10080) begin
        bht_bank_rd_data_out_1_142 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_142 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_143 <= 2'h0;
    end else if (bht_bank_sel_1_8_15) begin
      if (_T_10089) begin
        bht_bank_rd_data_out_1_143 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_143 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_144 <= 2'h0;
    end else if (bht_bank_sel_1_9_0) begin
      if (_T_10098) begin
        bht_bank_rd_data_out_1_144 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_144 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_145 <= 2'h0;
    end else if (bht_bank_sel_1_9_1) begin
      if (_T_10107) begin
        bht_bank_rd_data_out_1_145 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_145 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_146 <= 2'h0;
    end else if (bht_bank_sel_1_9_2) begin
      if (_T_10116) begin
        bht_bank_rd_data_out_1_146 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_146 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_147 <= 2'h0;
    end else if (bht_bank_sel_1_9_3) begin
      if (_T_10125) begin
        bht_bank_rd_data_out_1_147 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_147 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_148 <= 2'h0;
    end else if (bht_bank_sel_1_9_4) begin
      if (_T_10134) begin
        bht_bank_rd_data_out_1_148 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_148 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_149 <= 2'h0;
    end else if (bht_bank_sel_1_9_5) begin
      if (_T_10143) begin
        bht_bank_rd_data_out_1_149 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_149 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_150 <= 2'h0;
    end else if (bht_bank_sel_1_9_6) begin
      if (_T_10152) begin
        bht_bank_rd_data_out_1_150 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_150 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_151 <= 2'h0;
    end else if (bht_bank_sel_1_9_7) begin
      if (_T_10161) begin
        bht_bank_rd_data_out_1_151 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_151 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_152 <= 2'h0;
    end else if (bht_bank_sel_1_9_8) begin
      if (_T_10170) begin
        bht_bank_rd_data_out_1_152 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_152 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_153 <= 2'h0;
    end else if (bht_bank_sel_1_9_9) begin
      if (_T_10179) begin
        bht_bank_rd_data_out_1_153 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_153 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_154 <= 2'h0;
    end else if (bht_bank_sel_1_9_10) begin
      if (_T_10188) begin
        bht_bank_rd_data_out_1_154 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_154 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_155 <= 2'h0;
    end else if (bht_bank_sel_1_9_11) begin
      if (_T_10197) begin
        bht_bank_rd_data_out_1_155 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_155 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_156 <= 2'h0;
    end else if (bht_bank_sel_1_9_12) begin
      if (_T_10206) begin
        bht_bank_rd_data_out_1_156 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_156 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_157 <= 2'h0;
    end else if (bht_bank_sel_1_9_13) begin
      if (_T_10215) begin
        bht_bank_rd_data_out_1_157 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_157 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_158 <= 2'h0;
    end else if (bht_bank_sel_1_9_14) begin
      if (_T_10224) begin
        bht_bank_rd_data_out_1_158 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_158 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_159 <= 2'h0;
    end else if (bht_bank_sel_1_9_15) begin
      if (_T_10233) begin
        bht_bank_rd_data_out_1_159 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_159 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_160 <= 2'h0;
    end else if (bht_bank_sel_1_10_0) begin
      if (_T_10242) begin
        bht_bank_rd_data_out_1_160 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_160 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_161 <= 2'h0;
    end else if (bht_bank_sel_1_10_1) begin
      if (_T_10251) begin
        bht_bank_rd_data_out_1_161 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_161 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_162 <= 2'h0;
    end else if (bht_bank_sel_1_10_2) begin
      if (_T_10260) begin
        bht_bank_rd_data_out_1_162 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_162 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_163 <= 2'h0;
    end else if (bht_bank_sel_1_10_3) begin
      if (_T_10269) begin
        bht_bank_rd_data_out_1_163 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_163 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_164 <= 2'h0;
    end else if (bht_bank_sel_1_10_4) begin
      if (_T_10278) begin
        bht_bank_rd_data_out_1_164 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_164 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_165 <= 2'h0;
    end else if (bht_bank_sel_1_10_5) begin
      if (_T_10287) begin
        bht_bank_rd_data_out_1_165 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_165 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_166 <= 2'h0;
    end else if (bht_bank_sel_1_10_6) begin
      if (_T_10296) begin
        bht_bank_rd_data_out_1_166 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_166 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_167 <= 2'h0;
    end else if (bht_bank_sel_1_10_7) begin
      if (_T_10305) begin
        bht_bank_rd_data_out_1_167 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_167 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_168 <= 2'h0;
    end else if (bht_bank_sel_1_10_8) begin
      if (_T_10314) begin
        bht_bank_rd_data_out_1_168 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_168 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_169 <= 2'h0;
    end else if (bht_bank_sel_1_10_9) begin
      if (_T_10323) begin
        bht_bank_rd_data_out_1_169 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_169 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_170 <= 2'h0;
    end else if (bht_bank_sel_1_10_10) begin
      if (_T_10332) begin
        bht_bank_rd_data_out_1_170 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_170 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_171 <= 2'h0;
    end else if (bht_bank_sel_1_10_11) begin
      if (_T_10341) begin
        bht_bank_rd_data_out_1_171 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_171 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_172 <= 2'h0;
    end else if (bht_bank_sel_1_10_12) begin
      if (_T_10350) begin
        bht_bank_rd_data_out_1_172 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_172 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_173 <= 2'h0;
    end else if (bht_bank_sel_1_10_13) begin
      if (_T_10359) begin
        bht_bank_rd_data_out_1_173 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_173 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_174 <= 2'h0;
    end else if (bht_bank_sel_1_10_14) begin
      if (_T_10368) begin
        bht_bank_rd_data_out_1_174 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_174 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_175 <= 2'h0;
    end else if (bht_bank_sel_1_10_15) begin
      if (_T_10377) begin
        bht_bank_rd_data_out_1_175 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_175 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_176 <= 2'h0;
    end else if (bht_bank_sel_1_11_0) begin
      if (_T_10386) begin
        bht_bank_rd_data_out_1_176 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_176 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_177 <= 2'h0;
    end else if (bht_bank_sel_1_11_1) begin
      if (_T_10395) begin
        bht_bank_rd_data_out_1_177 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_177 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_178 <= 2'h0;
    end else if (bht_bank_sel_1_11_2) begin
      if (_T_10404) begin
        bht_bank_rd_data_out_1_178 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_178 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_179 <= 2'h0;
    end else if (bht_bank_sel_1_11_3) begin
      if (_T_10413) begin
        bht_bank_rd_data_out_1_179 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_179 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_180 <= 2'h0;
    end else if (bht_bank_sel_1_11_4) begin
      if (_T_10422) begin
        bht_bank_rd_data_out_1_180 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_180 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_181 <= 2'h0;
    end else if (bht_bank_sel_1_11_5) begin
      if (_T_10431) begin
        bht_bank_rd_data_out_1_181 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_181 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_182 <= 2'h0;
    end else if (bht_bank_sel_1_11_6) begin
      if (_T_10440) begin
        bht_bank_rd_data_out_1_182 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_182 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_183 <= 2'h0;
    end else if (bht_bank_sel_1_11_7) begin
      if (_T_10449) begin
        bht_bank_rd_data_out_1_183 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_183 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_184 <= 2'h0;
    end else if (bht_bank_sel_1_11_8) begin
      if (_T_10458) begin
        bht_bank_rd_data_out_1_184 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_184 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_185 <= 2'h0;
    end else if (bht_bank_sel_1_11_9) begin
      if (_T_10467) begin
        bht_bank_rd_data_out_1_185 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_185 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_186 <= 2'h0;
    end else if (bht_bank_sel_1_11_10) begin
      if (_T_10476) begin
        bht_bank_rd_data_out_1_186 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_186 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_187 <= 2'h0;
    end else if (bht_bank_sel_1_11_11) begin
      if (_T_10485) begin
        bht_bank_rd_data_out_1_187 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_187 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_188 <= 2'h0;
    end else if (bht_bank_sel_1_11_12) begin
      if (_T_10494) begin
        bht_bank_rd_data_out_1_188 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_188 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_189 <= 2'h0;
    end else if (bht_bank_sel_1_11_13) begin
      if (_T_10503) begin
        bht_bank_rd_data_out_1_189 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_189 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_190 <= 2'h0;
    end else if (bht_bank_sel_1_11_14) begin
      if (_T_10512) begin
        bht_bank_rd_data_out_1_190 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_190 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_191 <= 2'h0;
    end else if (bht_bank_sel_1_11_15) begin
      if (_T_10521) begin
        bht_bank_rd_data_out_1_191 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_191 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_192 <= 2'h0;
    end else if (bht_bank_sel_1_12_0) begin
      if (_T_10530) begin
        bht_bank_rd_data_out_1_192 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_192 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_193 <= 2'h0;
    end else if (bht_bank_sel_1_12_1) begin
      if (_T_10539) begin
        bht_bank_rd_data_out_1_193 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_193 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_194 <= 2'h0;
    end else if (bht_bank_sel_1_12_2) begin
      if (_T_10548) begin
        bht_bank_rd_data_out_1_194 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_194 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_195 <= 2'h0;
    end else if (bht_bank_sel_1_12_3) begin
      if (_T_10557) begin
        bht_bank_rd_data_out_1_195 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_195 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_196 <= 2'h0;
    end else if (bht_bank_sel_1_12_4) begin
      if (_T_10566) begin
        bht_bank_rd_data_out_1_196 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_196 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_197 <= 2'h0;
    end else if (bht_bank_sel_1_12_5) begin
      if (_T_10575) begin
        bht_bank_rd_data_out_1_197 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_197 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_198 <= 2'h0;
    end else if (bht_bank_sel_1_12_6) begin
      if (_T_10584) begin
        bht_bank_rd_data_out_1_198 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_198 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_199 <= 2'h0;
    end else if (bht_bank_sel_1_12_7) begin
      if (_T_10593) begin
        bht_bank_rd_data_out_1_199 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_199 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_200 <= 2'h0;
    end else if (bht_bank_sel_1_12_8) begin
      if (_T_10602) begin
        bht_bank_rd_data_out_1_200 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_200 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_201 <= 2'h0;
    end else if (bht_bank_sel_1_12_9) begin
      if (_T_10611) begin
        bht_bank_rd_data_out_1_201 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_201 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_202 <= 2'h0;
    end else if (bht_bank_sel_1_12_10) begin
      if (_T_10620) begin
        bht_bank_rd_data_out_1_202 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_202 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_203 <= 2'h0;
    end else if (bht_bank_sel_1_12_11) begin
      if (_T_10629) begin
        bht_bank_rd_data_out_1_203 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_203 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_204 <= 2'h0;
    end else if (bht_bank_sel_1_12_12) begin
      if (_T_10638) begin
        bht_bank_rd_data_out_1_204 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_204 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_205 <= 2'h0;
    end else if (bht_bank_sel_1_12_13) begin
      if (_T_10647) begin
        bht_bank_rd_data_out_1_205 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_205 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_206 <= 2'h0;
    end else if (bht_bank_sel_1_12_14) begin
      if (_T_10656) begin
        bht_bank_rd_data_out_1_206 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_206 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_207 <= 2'h0;
    end else if (bht_bank_sel_1_12_15) begin
      if (_T_10665) begin
        bht_bank_rd_data_out_1_207 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_207 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_208 <= 2'h0;
    end else if (bht_bank_sel_1_13_0) begin
      if (_T_10674) begin
        bht_bank_rd_data_out_1_208 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_208 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_209 <= 2'h0;
    end else if (bht_bank_sel_1_13_1) begin
      if (_T_10683) begin
        bht_bank_rd_data_out_1_209 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_209 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_210 <= 2'h0;
    end else if (bht_bank_sel_1_13_2) begin
      if (_T_10692) begin
        bht_bank_rd_data_out_1_210 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_210 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_211 <= 2'h0;
    end else if (bht_bank_sel_1_13_3) begin
      if (_T_10701) begin
        bht_bank_rd_data_out_1_211 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_211 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_212 <= 2'h0;
    end else if (bht_bank_sel_1_13_4) begin
      if (_T_10710) begin
        bht_bank_rd_data_out_1_212 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_212 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_213 <= 2'h0;
    end else if (bht_bank_sel_1_13_5) begin
      if (_T_10719) begin
        bht_bank_rd_data_out_1_213 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_213 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_214 <= 2'h0;
    end else if (bht_bank_sel_1_13_6) begin
      if (_T_10728) begin
        bht_bank_rd_data_out_1_214 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_214 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_215 <= 2'h0;
    end else if (bht_bank_sel_1_13_7) begin
      if (_T_10737) begin
        bht_bank_rd_data_out_1_215 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_215 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_216 <= 2'h0;
    end else if (bht_bank_sel_1_13_8) begin
      if (_T_10746) begin
        bht_bank_rd_data_out_1_216 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_216 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_217 <= 2'h0;
    end else if (bht_bank_sel_1_13_9) begin
      if (_T_10755) begin
        bht_bank_rd_data_out_1_217 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_217 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_218 <= 2'h0;
    end else if (bht_bank_sel_1_13_10) begin
      if (_T_10764) begin
        bht_bank_rd_data_out_1_218 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_218 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_219 <= 2'h0;
    end else if (bht_bank_sel_1_13_11) begin
      if (_T_10773) begin
        bht_bank_rd_data_out_1_219 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_219 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_220 <= 2'h0;
    end else if (bht_bank_sel_1_13_12) begin
      if (_T_10782) begin
        bht_bank_rd_data_out_1_220 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_220 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_221 <= 2'h0;
    end else if (bht_bank_sel_1_13_13) begin
      if (_T_10791) begin
        bht_bank_rd_data_out_1_221 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_221 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_222 <= 2'h0;
    end else if (bht_bank_sel_1_13_14) begin
      if (_T_10800) begin
        bht_bank_rd_data_out_1_222 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_222 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_223 <= 2'h0;
    end else if (bht_bank_sel_1_13_15) begin
      if (_T_10809) begin
        bht_bank_rd_data_out_1_223 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_223 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_224 <= 2'h0;
    end else if (bht_bank_sel_1_14_0) begin
      if (_T_10818) begin
        bht_bank_rd_data_out_1_224 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_224 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_225 <= 2'h0;
    end else if (bht_bank_sel_1_14_1) begin
      if (_T_10827) begin
        bht_bank_rd_data_out_1_225 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_225 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_226 <= 2'h0;
    end else if (bht_bank_sel_1_14_2) begin
      if (_T_10836) begin
        bht_bank_rd_data_out_1_226 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_226 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_227 <= 2'h0;
    end else if (bht_bank_sel_1_14_3) begin
      if (_T_10845) begin
        bht_bank_rd_data_out_1_227 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_227 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_228 <= 2'h0;
    end else if (bht_bank_sel_1_14_4) begin
      if (_T_10854) begin
        bht_bank_rd_data_out_1_228 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_228 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_229 <= 2'h0;
    end else if (bht_bank_sel_1_14_5) begin
      if (_T_10863) begin
        bht_bank_rd_data_out_1_229 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_229 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_230 <= 2'h0;
    end else if (bht_bank_sel_1_14_6) begin
      if (_T_10872) begin
        bht_bank_rd_data_out_1_230 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_230 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_231 <= 2'h0;
    end else if (bht_bank_sel_1_14_7) begin
      if (_T_10881) begin
        bht_bank_rd_data_out_1_231 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_231 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_232 <= 2'h0;
    end else if (bht_bank_sel_1_14_8) begin
      if (_T_10890) begin
        bht_bank_rd_data_out_1_232 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_232 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_233 <= 2'h0;
    end else if (bht_bank_sel_1_14_9) begin
      if (_T_10899) begin
        bht_bank_rd_data_out_1_233 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_233 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_234 <= 2'h0;
    end else if (bht_bank_sel_1_14_10) begin
      if (_T_10908) begin
        bht_bank_rd_data_out_1_234 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_234 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_235 <= 2'h0;
    end else if (bht_bank_sel_1_14_11) begin
      if (_T_10917) begin
        bht_bank_rd_data_out_1_235 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_235 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_236 <= 2'h0;
    end else if (bht_bank_sel_1_14_12) begin
      if (_T_10926) begin
        bht_bank_rd_data_out_1_236 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_236 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_237 <= 2'h0;
    end else if (bht_bank_sel_1_14_13) begin
      if (_T_10935) begin
        bht_bank_rd_data_out_1_237 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_237 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_238 <= 2'h0;
    end else if (bht_bank_sel_1_14_14) begin
      if (_T_10944) begin
        bht_bank_rd_data_out_1_238 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_238 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_239 <= 2'h0;
    end else if (bht_bank_sel_1_14_15) begin
      if (_T_10953) begin
        bht_bank_rd_data_out_1_239 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_239 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_240 <= 2'h0;
    end else if (bht_bank_sel_1_15_0) begin
      if (_T_10962) begin
        bht_bank_rd_data_out_1_240 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_240 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_241 <= 2'h0;
    end else if (bht_bank_sel_1_15_1) begin
      if (_T_10971) begin
        bht_bank_rd_data_out_1_241 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_241 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_242 <= 2'h0;
    end else if (bht_bank_sel_1_15_2) begin
      if (_T_10980) begin
        bht_bank_rd_data_out_1_242 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_242 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_243 <= 2'h0;
    end else if (bht_bank_sel_1_15_3) begin
      if (_T_10989) begin
        bht_bank_rd_data_out_1_243 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_243 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_244 <= 2'h0;
    end else if (bht_bank_sel_1_15_4) begin
      if (_T_10998) begin
        bht_bank_rd_data_out_1_244 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_244 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_245 <= 2'h0;
    end else if (bht_bank_sel_1_15_5) begin
      if (_T_11007) begin
        bht_bank_rd_data_out_1_245 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_245 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_246 <= 2'h0;
    end else if (bht_bank_sel_1_15_6) begin
      if (_T_11016) begin
        bht_bank_rd_data_out_1_246 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_246 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_247 <= 2'h0;
    end else if (bht_bank_sel_1_15_7) begin
      if (_T_11025) begin
        bht_bank_rd_data_out_1_247 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_247 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_248 <= 2'h0;
    end else if (bht_bank_sel_1_15_8) begin
      if (_T_11034) begin
        bht_bank_rd_data_out_1_248 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_248 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_249 <= 2'h0;
    end else if (bht_bank_sel_1_15_9) begin
      if (_T_11043) begin
        bht_bank_rd_data_out_1_249 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_249 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_250 <= 2'h0;
    end else if (bht_bank_sel_1_15_10) begin
      if (_T_11052) begin
        bht_bank_rd_data_out_1_250 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_250 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_251 <= 2'h0;
    end else if (bht_bank_sel_1_15_11) begin
      if (_T_11061) begin
        bht_bank_rd_data_out_1_251 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_251 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_252 <= 2'h0;
    end else if (bht_bank_sel_1_15_12) begin
      if (_T_11070) begin
        bht_bank_rd_data_out_1_252 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_252 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_253 <= 2'h0;
    end else if (bht_bank_sel_1_15_13) begin
      if (_T_11079) begin
        bht_bank_rd_data_out_1_253 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_253 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_254 <= 2'h0;
    end else if (bht_bank_sel_1_15_14) begin
      if (_T_11088) begin
        bht_bank_rd_data_out_1_254 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_254 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_255 <= 2'h0;
    end else if (bht_bank_sel_1_15_15) begin
      if (_T_11097) begin
        bht_bank_rd_data_out_1_255 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_255 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_0 <= 2'h0;
    end else if (bht_bank_sel_0_0_0) begin
      if (_T_6498) begin
        bht_bank_rd_data_out_0_0 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_0 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_1 <= 2'h0;
    end else if (bht_bank_sel_0_0_1) begin
      if (_T_6507) begin
        bht_bank_rd_data_out_0_1 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_1 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_2 <= 2'h0;
    end else if (bht_bank_sel_0_0_2) begin
      if (_T_6516) begin
        bht_bank_rd_data_out_0_2 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_2 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_3 <= 2'h0;
    end else if (bht_bank_sel_0_0_3) begin
      if (_T_6525) begin
        bht_bank_rd_data_out_0_3 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_3 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_4 <= 2'h0;
    end else if (bht_bank_sel_0_0_4) begin
      if (_T_6534) begin
        bht_bank_rd_data_out_0_4 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_4 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_5 <= 2'h0;
    end else if (bht_bank_sel_0_0_5) begin
      if (_T_6543) begin
        bht_bank_rd_data_out_0_5 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_5 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_6 <= 2'h0;
    end else if (bht_bank_sel_0_0_6) begin
      if (_T_6552) begin
        bht_bank_rd_data_out_0_6 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_6 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_7 <= 2'h0;
    end else if (bht_bank_sel_0_0_7) begin
      if (_T_6561) begin
        bht_bank_rd_data_out_0_7 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_7 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_8 <= 2'h0;
    end else if (bht_bank_sel_0_0_8) begin
      if (_T_6570) begin
        bht_bank_rd_data_out_0_8 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_8 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_9 <= 2'h0;
    end else if (bht_bank_sel_0_0_9) begin
      if (_T_6579) begin
        bht_bank_rd_data_out_0_9 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_9 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_10 <= 2'h0;
    end else if (bht_bank_sel_0_0_10) begin
      if (_T_6588) begin
        bht_bank_rd_data_out_0_10 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_10 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_11 <= 2'h0;
    end else if (bht_bank_sel_0_0_11) begin
      if (_T_6597) begin
        bht_bank_rd_data_out_0_11 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_11 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_12 <= 2'h0;
    end else if (bht_bank_sel_0_0_12) begin
      if (_T_6606) begin
        bht_bank_rd_data_out_0_12 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_12 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_13 <= 2'h0;
    end else if (bht_bank_sel_0_0_13) begin
      if (_T_6615) begin
        bht_bank_rd_data_out_0_13 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_13 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_14 <= 2'h0;
    end else if (bht_bank_sel_0_0_14) begin
      if (_T_6624) begin
        bht_bank_rd_data_out_0_14 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_14 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_15 <= 2'h0;
    end else if (bht_bank_sel_0_0_15) begin
      if (_T_6633) begin
        bht_bank_rd_data_out_0_15 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_15 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_16 <= 2'h0;
    end else if (bht_bank_sel_0_1_0) begin
      if (_T_6642) begin
        bht_bank_rd_data_out_0_16 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_16 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_17 <= 2'h0;
    end else if (bht_bank_sel_0_1_1) begin
      if (_T_6651) begin
        bht_bank_rd_data_out_0_17 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_17 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_18 <= 2'h0;
    end else if (bht_bank_sel_0_1_2) begin
      if (_T_6660) begin
        bht_bank_rd_data_out_0_18 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_18 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_19 <= 2'h0;
    end else if (bht_bank_sel_0_1_3) begin
      if (_T_6669) begin
        bht_bank_rd_data_out_0_19 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_19 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_20 <= 2'h0;
    end else if (bht_bank_sel_0_1_4) begin
      if (_T_6678) begin
        bht_bank_rd_data_out_0_20 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_20 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_21 <= 2'h0;
    end else if (bht_bank_sel_0_1_5) begin
      if (_T_6687) begin
        bht_bank_rd_data_out_0_21 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_21 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_22 <= 2'h0;
    end else if (bht_bank_sel_0_1_6) begin
      if (_T_6696) begin
        bht_bank_rd_data_out_0_22 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_22 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_23 <= 2'h0;
    end else if (bht_bank_sel_0_1_7) begin
      if (_T_6705) begin
        bht_bank_rd_data_out_0_23 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_23 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_24 <= 2'h0;
    end else if (bht_bank_sel_0_1_8) begin
      if (_T_6714) begin
        bht_bank_rd_data_out_0_24 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_24 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_25 <= 2'h0;
    end else if (bht_bank_sel_0_1_9) begin
      if (_T_6723) begin
        bht_bank_rd_data_out_0_25 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_25 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_26 <= 2'h0;
    end else if (bht_bank_sel_0_1_10) begin
      if (_T_6732) begin
        bht_bank_rd_data_out_0_26 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_26 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_27 <= 2'h0;
    end else if (bht_bank_sel_0_1_11) begin
      if (_T_6741) begin
        bht_bank_rd_data_out_0_27 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_27 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_28 <= 2'h0;
    end else if (bht_bank_sel_0_1_12) begin
      if (_T_6750) begin
        bht_bank_rd_data_out_0_28 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_28 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_29 <= 2'h0;
    end else if (bht_bank_sel_0_1_13) begin
      if (_T_6759) begin
        bht_bank_rd_data_out_0_29 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_29 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_30 <= 2'h0;
    end else if (bht_bank_sel_0_1_14) begin
      if (_T_6768) begin
        bht_bank_rd_data_out_0_30 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_30 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_31 <= 2'h0;
    end else if (bht_bank_sel_0_1_15) begin
      if (_T_6777) begin
        bht_bank_rd_data_out_0_31 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_31 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_32 <= 2'h0;
    end else if (bht_bank_sel_0_2_0) begin
      if (_T_6786) begin
        bht_bank_rd_data_out_0_32 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_32 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_33 <= 2'h0;
    end else if (bht_bank_sel_0_2_1) begin
      if (_T_6795) begin
        bht_bank_rd_data_out_0_33 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_33 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_34 <= 2'h0;
    end else if (bht_bank_sel_0_2_2) begin
      if (_T_6804) begin
        bht_bank_rd_data_out_0_34 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_34 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_35 <= 2'h0;
    end else if (bht_bank_sel_0_2_3) begin
      if (_T_6813) begin
        bht_bank_rd_data_out_0_35 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_35 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_36 <= 2'h0;
    end else if (bht_bank_sel_0_2_4) begin
      if (_T_6822) begin
        bht_bank_rd_data_out_0_36 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_36 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_37 <= 2'h0;
    end else if (bht_bank_sel_0_2_5) begin
      if (_T_6831) begin
        bht_bank_rd_data_out_0_37 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_37 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_38 <= 2'h0;
    end else if (bht_bank_sel_0_2_6) begin
      if (_T_6840) begin
        bht_bank_rd_data_out_0_38 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_38 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_39 <= 2'h0;
    end else if (bht_bank_sel_0_2_7) begin
      if (_T_6849) begin
        bht_bank_rd_data_out_0_39 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_39 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_40 <= 2'h0;
    end else if (bht_bank_sel_0_2_8) begin
      if (_T_6858) begin
        bht_bank_rd_data_out_0_40 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_40 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_41 <= 2'h0;
    end else if (bht_bank_sel_0_2_9) begin
      if (_T_6867) begin
        bht_bank_rd_data_out_0_41 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_41 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_42 <= 2'h0;
    end else if (bht_bank_sel_0_2_10) begin
      if (_T_6876) begin
        bht_bank_rd_data_out_0_42 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_42 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_43 <= 2'h0;
    end else if (bht_bank_sel_0_2_11) begin
      if (_T_6885) begin
        bht_bank_rd_data_out_0_43 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_43 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_44 <= 2'h0;
    end else if (bht_bank_sel_0_2_12) begin
      if (_T_6894) begin
        bht_bank_rd_data_out_0_44 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_44 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_45 <= 2'h0;
    end else if (bht_bank_sel_0_2_13) begin
      if (_T_6903) begin
        bht_bank_rd_data_out_0_45 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_45 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_46 <= 2'h0;
    end else if (bht_bank_sel_0_2_14) begin
      if (_T_6912) begin
        bht_bank_rd_data_out_0_46 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_46 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_47 <= 2'h0;
    end else if (bht_bank_sel_0_2_15) begin
      if (_T_6921) begin
        bht_bank_rd_data_out_0_47 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_47 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_48 <= 2'h0;
    end else if (bht_bank_sel_0_3_0) begin
      if (_T_6930) begin
        bht_bank_rd_data_out_0_48 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_48 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_49 <= 2'h0;
    end else if (bht_bank_sel_0_3_1) begin
      if (_T_6939) begin
        bht_bank_rd_data_out_0_49 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_49 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_50 <= 2'h0;
    end else if (bht_bank_sel_0_3_2) begin
      if (_T_6948) begin
        bht_bank_rd_data_out_0_50 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_50 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_51 <= 2'h0;
    end else if (bht_bank_sel_0_3_3) begin
      if (_T_6957) begin
        bht_bank_rd_data_out_0_51 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_51 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_52 <= 2'h0;
    end else if (bht_bank_sel_0_3_4) begin
      if (_T_6966) begin
        bht_bank_rd_data_out_0_52 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_52 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_53 <= 2'h0;
    end else if (bht_bank_sel_0_3_5) begin
      if (_T_6975) begin
        bht_bank_rd_data_out_0_53 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_53 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_54 <= 2'h0;
    end else if (bht_bank_sel_0_3_6) begin
      if (_T_6984) begin
        bht_bank_rd_data_out_0_54 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_54 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_55 <= 2'h0;
    end else if (bht_bank_sel_0_3_7) begin
      if (_T_6993) begin
        bht_bank_rd_data_out_0_55 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_55 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_56 <= 2'h0;
    end else if (bht_bank_sel_0_3_8) begin
      if (_T_7002) begin
        bht_bank_rd_data_out_0_56 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_56 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_57 <= 2'h0;
    end else if (bht_bank_sel_0_3_9) begin
      if (_T_7011) begin
        bht_bank_rd_data_out_0_57 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_57 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_58 <= 2'h0;
    end else if (bht_bank_sel_0_3_10) begin
      if (_T_7020) begin
        bht_bank_rd_data_out_0_58 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_58 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_59 <= 2'h0;
    end else if (bht_bank_sel_0_3_11) begin
      if (_T_7029) begin
        bht_bank_rd_data_out_0_59 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_59 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_60 <= 2'h0;
    end else if (bht_bank_sel_0_3_12) begin
      if (_T_7038) begin
        bht_bank_rd_data_out_0_60 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_60 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_61 <= 2'h0;
    end else if (bht_bank_sel_0_3_13) begin
      if (_T_7047) begin
        bht_bank_rd_data_out_0_61 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_61 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_62 <= 2'h0;
    end else if (bht_bank_sel_0_3_14) begin
      if (_T_7056) begin
        bht_bank_rd_data_out_0_62 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_62 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_63 <= 2'h0;
    end else if (bht_bank_sel_0_3_15) begin
      if (_T_7065) begin
        bht_bank_rd_data_out_0_63 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_63 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_64 <= 2'h0;
    end else if (bht_bank_sel_0_4_0) begin
      if (_T_7074) begin
        bht_bank_rd_data_out_0_64 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_64 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_65 <= 2'h0;
    end else if (bht_bank_sel_0_4_1) begin
      if (_T_7083) begin
        bht_bank_rd_data_out_0_65 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_65 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_66 <= 2'h0;
    end else if (bht_bank_sel_0_4_2) begin
      if (_T_7092) begin
        bht_bank_rd_data_out_0_66 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_66 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_67 <= 2'h0;
    end else if (bht_bank_sel_0_4_3) begin
      if (_T_7101) begin
        bht_bank_rd_data_out_0_67 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_67 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_68 <= 2'h0;
    end else if (bht_bank_sel_0_4_4) begin
      if (_T_7110) begin
        bht_bank_rd_data_out_0_68 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_68 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_69 <= 2'h0;
    end else if (bht_bank_sel_0_4_5) begin
      if (_T_7119) begin
        bht_bank_rd_data_out_0_69 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_69 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_70 <= 2'h0;
    end else if (bht_bank_sel_0_4_6) begin
      if (_T_7128) begin
        bht_bank_rd_data_out_0_70 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_70 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_71 <= 2'h0;
    end else if (bht_bank_sel_0_4_7) begin
      if (_T_7137) begin
        bht_bank_rd_data_out_0_71 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_71 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_72 <= 2'h0;
    end else if (bht_bank_sel_0_4_8) begin
      if (_T_7146) begin
        bht_bank_rd_data_out_0_72 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_72 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_73 <= 2'h0;
    end else if (bht_bank_sel_0_4_9) begin
      if (_T_7155) begin
        bht_bank_rd_data_out_0_73 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_73 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_74 <= 2'h0;
    end else if (bht_bank_sel_0_4_10) begin
      if (_T_7164) begin
        bht_bank_rd_data_out_0_74 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_74 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_75 <= 2'h0;
    end else if (bht_bank_sel_0_4_11) begin
      if (_T_7173) begin
        bht_bank_rd_data_out_0_75 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_75 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_76 <= 2'h0;
    end else if (bht_bank_sel_0_4_12) begin
      if (_T_7182) begin
        bht_bank_rd_data_out_0_76 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_76 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_77 <= 2'h0;
    end else if (bht_bank_sel_0_4_13) begin
      if (_T_7191) begin
        bht_bank_rd_data_out_0_77 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_77 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_78 <= 2'h0;
    end else if (bht_bank_sel_0_4_14) begin
      if (_T_7200) begin
        bht_bank_rd_data_out_0_78 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_78 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_79 <= 2'h0;
    end else if (bht_bank_sel_0_4_15) begin
      if (_T_7209) begin
        bht_bank_rd_data_out_0_79 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_79 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_80 <= 2'h0;
    end else if (bht_bank_sel_0_5_0) begin
      if (_T_7218) begin
        bht_bank_rd_data_out_0_80 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_80 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_81 <= 2'h0;
    end else if (bht_bank_sel_0_5_1) begin
      if (_T_7227) begin
        bht_bank_rd_data_out_0_81 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_81 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_82 <= 2'h0;
    end else if (bht_bank_sel_0_5_2) begin
      if (_T_7236) begin
        bht_bank_rd_data_out_0_82 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_82 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_83 <= 2'h0;
    end else if (bht_bank_sel_0_5_3) begin
      if (_T_7245) begin
        bht_bank_rd_data_out_0_83 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_83 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_84 <= 2'h0;
    end else if (bht_bank_sel_0_5_4) begin
      if (_T_7254) begin
        bht_bank_rd_data_out_0_84 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_84 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_85 <= 2'h0;
    end else if (bht_bank_sel_0_5_5) begin
      if (_T_7263) begin
        bht_bank_rd_data_out_0_85 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_85 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_86 <= 2'h0;
    end else if (bht_bank_sel_0_5_6) begin
      if (_T_7272) begin
        bht_bank_rd_data_out_0_86 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_86 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_87 <= 2'h0;
    end else if (bht_bank_sel_0_5_7) begin
      if (_T_7281) begin
        bht_bank_rd_data_out_0_87 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_87 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_88 <= 2'h0;
    end else if (bht_bank_sel_0_5_8) begin
      if (_T_7290) begin
        bht_bank_rd_data_out_0_88 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_88 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_89 <= 2'h0;
    end else if (bht_bank_sel_0_5_9) begin
      if (_T_7299) begin
        bht_bank_rd_data_out_0_89 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_89 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_90 <= 2'h0;
    end else if (bht_bank_sel_0_5_10) begin
      if (_T_7308) begin
        bht_bank_rd_data_out_0_90 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_90 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_91 <= 2'h0;
    end else if (bht_bank_sel_0_5_11) begin
      if (_T_7317) begin
        bht_bank_rd_data_out_0_91 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_91 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_92 <= 2'h0;
    end else if (bht_bank_sel_0_5_12) begin
      if (_T_7326) begin
        bht_bank_rd_data_out_0_92 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_92 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_93 <= 2'h0;
    end else if (bht_bank_sel_0_5_13) begin
      if (_T_7335) begin
        bht_bank_rd_data_out_0_93 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_93 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_94 <= 2'h0;
    end else if (bht_bank_sel_0_5_14) begin
      if (_T_7344) begin
        bht_bank_rd_data_out_0_94 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_94 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_95 <= 2'h0;
    end else if (bht_bank_sel_0_5_15) begin
      if (_T_7353) begin
        bht_bank_rd_data_out_0_95 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_95 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_96 <= 2'h0;
    end else if (bht_bank_sel_0_6_0) begin
      if (_T_7362) begin
        bht_bank_rd_data_out_0_96 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_96 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_97 <= 2'h0;
    end else if (bht_bank_sel_0_6_1) begin
      if (_T_7371) begin
        bht_bank_rd_data_out_0_97 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_97 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_98 <= 2'h0;
    end else if (bht_bank_sel_0_6_2) begin
      if (_T_7380) begin
        bht_bank_rd_data_out_0_98 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_98 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_99 <= 2'h0;
    end else if (bht_bank_sel_0_6_3) begin
      if (_T_7389) begin
        bht_bank_rd_data_out_0_99 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_99 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_100 <= 2'h0;
    end else if (bht_bank_sel_0_6_4) begin
      if (_T_7398) begin
        bht_bank_rd_data_out_0_100 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_100 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_101 <= 2'h0;
    end else if (bht_bank_sel_0_6_5) begin
      if (_T_7407) begin
        bht_bank_rd_data_out_0_101 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_101 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_102 <= 2'h0;
    end else if (bht_bank_sel_0_6_6) begin
      if (_T_7416) begin
        bht_bank_rd_data_out_0_102 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_102 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_103 <= 2'h0;
    end else if (bht_bank_sel_0_6_7) begin
      if (_T_7425) begin
        bht_bank_rd_data_out_0_103 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_103 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_104 <= 2'h0;
    end else if (bht_bank_sel_0_6_8) begin
      if (_T_7434) begin
        bht_bank_rd_data_out_0_104 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_104 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_105 <= 2'h0;
    end else if (bht_bank_sel_0_6_9) begin
      if (_T_7443) begin
        bht_bank_rd_data_out_0_105 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_105 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_106 <= 2'h0;
    end else if (bht_bank_sel_0_6_10) begin
      if (_T_7452) begin
        bht_bank_rd_data_out_0_106 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_106 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_107 <= 2'h0;
    end else if (bht_bank_sel_0_6_11) begin
      if (_T_7461) begin
        bht_bank_rd_data_out_0_107 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_107 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_108 <= 2'h0;
    end else if (bht_bank_sel_0_6_12) begin
      if (_T_7470) begin
        bht_bank_rd_data_out_0_108 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_108 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_109 <= 2'h0;
    end else if (bht_bank_sel_0_6_13) begin
      if (_T_7479) begin
        bht_bank_rd_data_out_0_109 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_109 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_110 <= 2'h0;
    end else if (bht_bank_sel_0_6_14) begin
      if (_T_7488) begin
        bht_bank_rd_data_out_0_110 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_110 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_111 <= 2'h0;
    end else if (bht_bank_sel_0_6_15) begin
      if (_T_7497) begin
        bht_bank_rd_data_out_0_111 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_111 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_112 <= 2'h0;
    end else if (bht_bank_sel_0_7_0) begin
      if (_T_7506) begin
        bht_bank_rd_data_out_0_112 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_112 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_113 <= 2'h0;
    end else if (bht_bank_sel_0_7_1) begin
      if (_T_7515) begin
        bht_bank_rd_data_out_0_113 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_113 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_114 <= 2'h0;
    end else if (bht_bank_sel_0_7_2) begin
      if (_T_7524) begin
        bht_bank_rd_data_out_0_114 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_114 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_115 <= 2'h0;
    end else if (bht_bank_sel_0_7_3) begin
      if (_T_7533) begin
        bht_bank_rd_data_out_0_115 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_115 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_116 <= 2'h0;
    end else if (bht_bank_sel_0_7_4) begin
      if (_T_7542) begin
        bht_bank_rd_data_out_0_116 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_116 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_117 <= 2'h0;
    end else if (bht_bank_sel_0_7_5) begin
      if (_T_7551) begin
        bht_bank_rd_data_out_0_117 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_117 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_118 <= 2'h0;
    end else if (bht_bank_sel_0_7_6) begin
      if (_T_7560) begin
        bht_bank_rd_data_out_0_118 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_118 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_119 <= 2'h0;
    end else if (bht_bank_sel_0_7_7) begin
      if (_T_7569) begin
        bht_bank_rd_data_out_0_119 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_119 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_120 <= 2'h0;
    end else if (bht_bank_sel_0_7_8) begin
      if (_T_7578) begin
        bht_bank_rd_data_out_0_120 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_120 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_121 <= 2'h0;
    end else if (bht_bank_sel_0_7_9) begin
      if (_T_7587) begin
        bht_bank_rd_data_out_0_121 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_121 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_122 <= 2'h0;
    end else if (bht_bank_sel_0_7_10) begin
      if (_T_7596) begin
        bht_bank_rd_data_out_0_122 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_122 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_123 <= 2'h0;
    end else if (bht_bank_sel_0_7_11) begin
      if (_T_7605) begin
        bht_bank_rd_data_out_0_123 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_123 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_124 <= 2'h0;
    end else if (bht_bank_sel_0_7_12) begin
      if (_T_7614) begin
        bht_bank_rd_data_out_0_124 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_124 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_125 <= 2'h0;
    end else if (bht_bank_sel_0_7_13) begin
      if (_T_7623) begin
        bht_bank_rd_data_out_0_125 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_125 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_126 <= 2'h0;
    end else if (bht_bank_sel_0_7_14) begin
      if (_T_7632) begin
        bht_bank_rd_data_out_0_126 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_126 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_127 <= 2'h0;
    end else if (bht_bank_sel_0_7_15) begin
      if (_T_7641) begin
        bht_bank_rd_data_out_0_127 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_127 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_128 <= 2'h0;
    end else if (bht_bank_sel_0_8_0) begin
      if (_T_7650) begin
        bht_bank_rd_data_out_0_128 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_128 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_129 <= 2'h0;
    end else if (bht_bank_sel_0_8_1) begin
      if (_T_7659) begin
        bht_bank_rd_data_out_0_129 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_129 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_130 <= 2'h0;
    end else if (bht_bank_sel_0_8_2) begin
      if (_T_7668) begin
        bht_bank_rd_data_out_0_130 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_130 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_131 <= 2'h0;
    end else if (bht_bank_sel_0_8_3) begin
      if (_T_7677) begin
        bht_bank_rd_data_out_0_131 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_131 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_132 <= 2'h0;
    end else if (bht_bank_sel_0_8_4) begin
      if (_T_7686) begin
        bht_bank_rd_data_out_0_132 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_132 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_133 <= 2'h0;
    end else if (bht_bank_sel_0_8_5) begin
      if (_T_7695) begin
        bht_bank_rd_data_out_0_133 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_133 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_134 <= 2'h0;
    end else if (bht_bank_sel_0_8_6) begin
      if (_T_7704) begin
        bht_bank_rd_data_out_0_134 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_134 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_135 <= 2'h0;
    end else if (bht_bank_sel_0_8_7) begin
      if (_T_7713) begin
        bht_bank_rd_data_out_0_135 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_135 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_136 <= 2'h0;
    end else if (bht_bank_sel_0_8_8) begin
      if (_T_7722) begin
        bht_bank_rd_data_out_0_136 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_136 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_137 <= 2'h0;
    end else if (bht_bank_sel_0_8_9) begin
      if (_T_7731) begin
        bht_bank_rd_data_out_0_137 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_137 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_138 <= 2'h0;
    end else if (bht_bank_sel_0_8_10) begin
      if (_T_7740) begin
        bht_bank_rd_data_out_0_138 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_138 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_139 <= 2'h0;
    end else if (bht_bank_sel_0_8_11) begin
      if (_T_7749) begin
        bht_bank_rd_data_out_0_139 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_139 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_140 <= 2'h0;
    end else if (bht_bank_sel_0_8_12) begin
      if (_T_7758) begin
        bht_bank_rd_data_out_0_140 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_140 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_141 <= 2'h0;
    end else if (bht_bank_sel_0_8_13) begin
      if (_T_7767) begin
        bht_bank_rd_data_out_0_141 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_141 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_142 <= 2'h0;
    end else if (bht_bank_sel_0_8_14) begin
      if (_T_7776) begin
        bht_bank_rd_data_out_0_142 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_142 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_143 <= 2'h0;
    end else if (bht_bank_sel_0_8_15) begin
      if (_T_7785) begin
        bht_bank_rd_data_out_0_143 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_143 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_144 <= 2'h0;
    end else if (bht_bank_sel_0_9_0) begin
      if (_T_7794) begin
        bht_bank_rd_data_out_0_144 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_144 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_145 <= 2'h0;
    end else if (bht_bank_sel_0_9_1) begin
      if (_T_7803) begin
        bht_bank_rd_data_out_0_145 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_145 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_146 <= 2'h0;
    end else if (bht_bank_sel_0_9_2) begin
      if (_T_7812) begin
        bht_bank_rd_data_out_0_146 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_146 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_147 <= 2'h0;
    end else if (bht_bank_sel_0_9_3) begin
      if (_T_7821) begin
        bht_bank_rd_data_out_0_147 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_147 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_148 <= 2'h0;
    end else if (bht_bank_sel_0_9_4) begin
      if (_T_7830) begin
        bht_bank_rd_data_out_0_148 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_148 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_149 <= 2'h0;
    end else if (bht_bank_sel_0_9_5) begin
      if (_T_7839) begin
        bht_bank_rd_data_out_0_149 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_149 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_150 <= 2'h0;
    end else if (bht_bank_sel_0_9_6) begin
      if (_T_7848) begin
        bht_bank_rd_data_out_0_150 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_150 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_151 <= 2'h0;
    end else if (bht_bank_sel_0_9_7) begin
      if (_T_7857) begin
        bht_bank_rd_data_out_0_151 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_151 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_152 <= 2'h0;
    end else if (bht_bank_sel_0_9_8) begin
      if (_T_7866) begin
        bht_bank_rd_data_out_0_152 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_152 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_153 <= 2'h0;
    end else if (bht_bank_sel_0_9_9) begin
      if (_T_7875) begin
        bht_bank_rd_data_out_0_153 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_153 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_154 <= 2'h0;
    end else if (bht_bank_sel_0_9_10) begin
      if (_T_7884) begin
        bht_bank_rd_data_out_0_154 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_154 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_155 <= 2'h0;
    end else if (bht_bank_sel_0_9_11) begin
      if (_T_7893) begin
        bht_bank_rd_data_out_0_155 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_155 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_156 <= 2'h0;
    end else if (bht_bank_sel_0_9_12) begin
      if (_T_7902) begin
        bht_bank_rd_data_out_0_156 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_156 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_157 <= 2'h0;
    end else if (bht_bank_sel_0_9_13) begin
      if (_T_7911) begin
        bht_bank_rd_data_out_0_157 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_157 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_158 <= 2'h0;
    end else if (bht_bank_sel_0_9_14) begin
      if (_T_7920) begin
        bht_bank_rd_data_out_0_158 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_158 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_159 <= 2'h0;
    end else if (bht_bank_sel_0_9_15) begin
      if (_T_7929) begin
        bht_bank_rd_data_out_0_159 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_159 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_160 <= 2'h0;
    end else if (bht_bank_sel_0_10_0) begin
      if (_T_7938) begin
        bht_bank_rd_data_out_0_160 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_160 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_161 <= 2'h0;
    end else if (bht_bank_sel_0_10_1) begin
      if (_T_7947) begin
        bht_bank_rd_data_out_0_161 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_161 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_162 <= 2'h0;
    end else if (bht_bank_sel_0_10_2) begin
      if (_T_7956) begin
        bht_bank_rd_data_out_0_162 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_162 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_163 <= 2'h0;
    end else if (bht_bank_sel_0_10_3) begin
      if (_T_7965) begin
        bht_bank_rd_data_out_0_163 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_163 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_164 <= 2'h0;
    end else if (bht_bank_sel_0_10_4) begin
      if (_T_7974) begin
        bht_bank_rd_data_out_0_164 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_164 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_165 <= 2'h0;
    end else if (bht_bank_sel_0_10_5) begin
      if (_T_7983) begin
        bht_bank_rd_data_out_0_165 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_165 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_166 <= 2'h0;
    end else if (bht_bank_sel_0_10_6) begin
      if (_T_7992) begin
        bht_bank_rd_data_out_0_166 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_166 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_167 <= 2'h0;
    end else if (bht_bank_sel_0_10_7) begin
      if (_T_8001) begin
        bht_bank_rd_data_out_0_167 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_167 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_168 <= 2'h0;
    end else if (bht_bank_sel_0_10_8) begin
      if (_T_8010) begin
        bht_bank_rd_data_out_0_168 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_168 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_169 <= 2'h0;
    end else if (bht_bank_sel_0_10_9) begin
      if (_T_8019) begin
        bht_bank_rd_data_out_0_169 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_169 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_170 <= 2'h0;
    end else if (bht_bank_sel_0_10_10) begin
      if (_T_8028) begin
        bht_bank_rd_data_out_0_170 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_170 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_171 <= 2'h0;
    end else if (bht_bank_sel_0_10_11) begin
      if (_T_8037) begin
        bht_bank_rd_data_out_0_171 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_171 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_172 <= 2'h0;
    end else if (bht_bank_sel_0_10_12) begin
      if (_T_8046) begin
        bht_bank_rd_data_out_0_172 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_172 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_173 <= 2'h0;
    end else if (bht_bank_sel_0_10_13) begin
      if (_T_8055) begin
        bht_bank_rd_data_out_0_173 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_173 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_174 <= 2'h0;
    end else if (bht_bank_sel_0_10_14) begin
      if (_T_8064) begin
        bht_bank_rd_data_out_0_174 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_174 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_175 <= 2'h0;
    end else if (bht_bank_sel_0_10_15) begin
      if (_T_8073) begin
        bht_bank_rd_data_out_0_175 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_175 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_176 <= 2'h0;
    end else if (bht_bank_sel_0_11_0) begin
      if (_T_8082) begin
        bht_bank_rd_data_out_0_176 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_176 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_177 <= 2'h0;
    end else if (bht_bank_sel_0_11_1) begin
      if (_T_8091) begin
        bht_bank_rd_data_out_0_177 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_177 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_178 <= 2'h0;
    end else if (bht_bank_sel_0_11_2) begin
      if (_T_8100) begin
        bht_bank_rd_data_out_0_178 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_178 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_179 <= 2'h0;
    end else if (bht_bank_sel_0_11_3) begin
      if (_T_8109) begin
        bht_bank_rd_data_out_0_179 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_179 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_180 <= 2'h0;
    end else if (bht_bank_sel_0_11_4) begin
      if (_T_8118) begin
        bht_bank_rd_data_out_0_180 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_180 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_181 <= 2'h0;
    end else if (bht_bank_sel_0_11_5) begin
      if (_T_8127) begin
        bht_bank_rd_data_out_0_181 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_181 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_182 <= 2'h0;
    end else if (bht_bank_sel_0_11_6) begin
      if (_T_8136) begin
        bht_bank_rd_data_out_0_182 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_182 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_183 <= 2'h0;
    end else if (bht_bank_sel_0_11_7) begin
      if (_T_8145) begin
        bht_bank_rd_data_out_0_183 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_183 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_184 <= 2'h0;
    end else if (bht_bank_sel_0_11_8) begin
      if (_T_8154) begin
        bht_bank_rd_data_out_0_184 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_184 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_185 <= 2'h0;
    end else if (bht_bank_sel_0_11_9) begin
      if (_T_8163) begin
        bht_bank_rd_data_out_0_185 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_185 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_186 <= 2'h0;
    end else if (bht_bank_sel_0_11_10) begin
      if (_T_8172) begin
        bht_bank_rd_data_out_0_186 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_186 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_187 <= 2'h0;
    end else if (bht_bank_sel_0_11_11) begin
      if (_T_8181) begin
        bht_bank_rd_data_out_0_187 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_187 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_188 <= 2'h0;
    end else if (bht_bank_sel_0_11_12) begin
      if (_T_8190) begin
        bht_bank_rd_data_out_0_188 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_188 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_189 <= 2'h0;
    end else if (bht_bank_sel_0_11_13) begin
      if (_T_8199) begin
        bht_bank_rd_data_out_0_189 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_189 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_190 <= 2'h0;
    end else if (bht_bank_sel_0_11_14) begin
      if (_T_8208) begin
        bht_bank_rd_data_out_0_190 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_190 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_191 <= 2'h0;
    end else if (bht_bank_sel_0_11_15) begin
      if (_T_8217) begin
        bht_bank_rd_data_out_0_191 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_191 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_192 <= 2'h0;
    end else if (bht_bank_sel_0_12_0) begin
      if (_T_8226) begin
        bht_bank_rd_data_out_0_192 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_192 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_193 <= 2'h0;
    end else if (bht_bank_sel_0_12_1) begin
      if (_T_8235) begin
        bht_bank_rd_data_out_0_193 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_193 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_194 <= 2'h0;
    end else if (bht_bank_sel_0_12_2) begin
      if (_T_8244) begin
        bht_bank_rd_data_out_0_194 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_194 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_195 <= 2'h0;
    end else if (bht_bank_sel_0_12_3) begin
      if (_T_8253) begin
        bht_bank_rd_data_out_0_195 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_195 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_196 <= 2'h0;
    end else if (bht_bank_sel_0_12_4) begin
      if (_T_8262) begin
        bht_bank_rd_data_out_0_196 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_196 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_197 <= 2'h0;
    end else if (bht_bank_sel_0_12_5) begin
      if (_T_8271) begin
        bht_bank_rd_data_out_0_197 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_197 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_198 <= 2'h0;
    end else if (bht_bank_sel_0_12_6) begin
      if (_T_8280) begin
        bht_bank_rd_data_out_0_198 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_198 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_199 <= 2'h0;
    end else if (bht_bank_sel_0_12_7) begin
      if (_T_8289) begin
        bht_bank_rd_data_out_0_199 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_199 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_200 <= 2'h0;
    end else if (bht_bank_sel_0_12_8) begin
      if (_T_8298) begin
        bht_bank_rd_data_out_0_200 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_200 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_201 <= 2'h0;
    end else if (bht_bank_sel_0_12_9) begin
      if (_T_8307) begin
        bht_bank_rd_data_out_0_201 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_201 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_202 <= 2'h0;
    end else if (bht_bank_sel_0_12_10) begin
      if (_T_8316) begin
        bht_bank_rd_data_out_0_202 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_202 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_203 <= 2'h0;
    end else if (bht_bank_sel_0_12_11) begin
      if (_T_8325) begin
        bht_bank_rd_data_out_0_203 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_203 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_204 <= 2'h0;
    end else if (bht_bank_sel_0_12_12) begin
      if (_T_8334) begin
        bht_bank_rd_data_out_0_204 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_204 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_205 <= 2'h0;
    end else if (bht_bank_sel_0_12_13) begin
      if (_T_8343) begin
        bht_bank_rd_data_out_0_205 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_205 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_206 <= 2'h0;
    end else if (bht_bank_sel_0_12_14) begin
      if (_T_8352) begin
        bht_bank_rd_data_out_0_206 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_206 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_207 <= 2'h0;
    end else if (bht_bank_sel_0_12_15) begin
      if (_T_8361) begin
        bht_bank_rd_data_out_0_207 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_207 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_208 <= 2'h0;
    end else if (bht_bank_sel_0_13_0) begin
      if (_T_8370) begin
        bht_bank_rd_data_out_0_208 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_208 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_209 <= 2'h0;
    end else if (bht_bank_sel_0_13_1) begin
      if (_T_8379) begin
        bht_bank_rd_data_out_0_209 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_209 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_210 <= 2'h0;
    end else if (bht_bank_sel_0_13_2) begin
      if (_T_8388) begin
        bht_bank_rd_data_out_0_210 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_210 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_211 <= 2'h0;
    end else if (bht_bank_sel_0_13_3) begin
      if (_T_8397) begin
        bht_bank_rd_data_out_0_211 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_211 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_212 <= 2'h0;
    end else if (bht_bank_sel_0_13_4) begin
      if (_T_8406) begin
        bht_bank_rd_data_out_0_212 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_212 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_213 <= 2'h0;
    end else if (bht_bank_sel_0_13_5) begin
      if (_T_8415) begin
        bht_bank_rd_data_out_0_213 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_213 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_214 <= 2'h0;
    end else if (bht_bank_sel_0_13_6) begin
      if (_T_8424) begin
        bht_bank_rd_data_out_0_214 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_214 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_215 <= 2'h0;
    end else if (bht_bank_sel_0_13_7) begin
      if (_T_8433) begin
        bht_bank_rd_data_out_0_215 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_215 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_216 <= 2'h0;
    end else if (bht_bank_sel_0_13_8) begin
      if (_T_8442) begin
        bht_bank_rd_data_out_0_216 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_216 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_217 <= 2'h0;
    end else if (bht_bank_sel_0_13_9) begin
      if (_T_8451) begin
        bht_bank_rd_data_out_0_217 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_217 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_218 <= 2'h0;
    end else if (bht_bank_sel_0_13_10) begin
      if (_T_8460) begin
        bht_bank_rd_data_out_0_218 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_218 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_219 <= 2'h0;
    end else if (bht_bank_sel_0_13_11) begin
      if (_T_8469) begin
        bht_bank_rd_data_out_0_219 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_219 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_220 <= 2'h0;
    end else if (bht_bank_sel_0_13_12) begin
      if (_T_8478) begin
        bht_bank_rd_data_out_0_220 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_220 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_221 <= 2'h0;
    end else if (bht_bank_sel_0_13_13) begin
      if (_T_8487) begin
        bht_bank_rd_data_out_0_221 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_221 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_222 <= 2'h0;
    end else if (bht_bank_sel_0_13_14) begin
      if (_T_8496) begin
        bht_bank_rd_data_out_0_222 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_222 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_223 <= 2'h0;
    end else if (bht_bank_sel_0_13_15) begin
      if (_T_8505) begin
        bht_bank_rd_data_out_0_223 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_223 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_224 <= 2'h0;
    end else if (bht_bank_sel_0_14_0) begin
      if (_T_8514) begin
        bht_bank_rd_data_out_0_224 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_224 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_225 <= 2'h0;
    end else if (bht_bank_sel_0_14_1) begin
      if (_T_8523) begin
        bht_bank_rd_data_out_0_225 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_225 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_226 <= 2'h0;
    end else if (bht_bank_sel_0_14_2) begin
      if (_T_8532) begin
        bht_bank_rd_data_out_0_226 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_226 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_227 <= 2'h0;
    end else if (bht_bank_sel_0_14_3) begin
      if (_T_8541) begin
        bht_bank_rd_data_out_0_227 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_227 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_228 <= 2'h0;
    end else if (bht_bank_sel_0_14_4) begin
      if (_T_8550) begin
        bht_bank_rd_data_out_0_228 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_228 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_229 <= 2'h0;
    end else if (bht_bank_sel_0_14_5) begin
      if (_T_8559) begin
        bht_bank_rd_data_out_0_229 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_229 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_230 <= 2'h0;
    end else if (bht_bank_sel_0_14_6) begin
      if (_T_8568) begin
        bht_bank_rd_data_out_0_230 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_230 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_231 <= 2'h0;
    end else if (bht_bank_sel_0_14_7) begin
      if (_T_8577) begin
        bht_bank_rd_data_out_0_231 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_231 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_232 <= 2'h0;
    end else if (bht_bank_sel_0_14_8) begin
      if (_T_8586) begin
        bht_bank_rd_data_out_0_232 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_232 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_233 <= 2'h0;
    end else if (bht_bank_sel_0_14_9) begin
      if (_T_8595) begin
        bht_bank_rd_data_out_0_233 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_233 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_234 <= 2'h0;
    end else if (bht_bank_sel_0_14_10) begin
      if (_T_8604) begin
        bht_bank_rd_data_out_0_234 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_234 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_235 <= 2'h0;
    end else if (bht_bank_sel_0_14_11) begin
      if (_T_8613) begin
        bht_bank_rd_data_out_0_235 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_235 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_236 <= 2'h0;
    end else if (bht_bank_sel_0_14_12) begin
      if (_T_8622) begin
        bht_bank_rd_data_out_0_236 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_236 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_237 <= 2'h0;
    end else if (bht_bank_sel_0_14_13) begin
      if (_T_8631) begin
        bht_bank_rd_data_out_0_237 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_237 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_238 <= 2'h0;
    end else if (bht_bank_sel_0_14_14) begin
      if (_T_8640) begin
        bht_bank_rd_data_out_0_238 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_238 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_239 <= 2'h0;
    end else if (bht_bank_sel_0_14_15) begin
      if (_T_8649) begin
        bht_bank_rd_data_out_0_239 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_239 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_240 <= 2'h0;
    end else if (bht_bank_sel_0_15_0) begin
      if (_T_8658) begin
        bht_bank_rd_data_out_0_240 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_240 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_241 <= 2'h0;
    end else if (bht_bank_sel_0_15_1) begin
      if (_T_8667) begin
        bht_bank_rd_data_out_0_241 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_241 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_242 <= 2'h0;
    end else if (bht_bank_sel_0_15_2) begin
      if (_T_8676) begin
        bht_bank_rd_data_out_0_242 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_242 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_243 <= 2'h0;
    end else if (bht_bank_sel_0_15_3) begin
      if (_T_8685) begin
        bht_bank_rd_data_out_0_243 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_243 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_244 <= 2'h0;
    end else if (bht_bank_sel_0_15_4) begin
      if (_T_8694) begin
        bht_bank_rd_data_out_0_244 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_244 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_245 <= 2'h0;
    end else if (bht_bank_sel_0_15_5) begin
      if (_T_8703) begin
        bht_bank_rd_data_out_0_245 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_245 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_246 <= 2'h0;
    end else if (bht_bank_sel_0_15_6) begin
      if (_T_8712) begin
        bht_bank_rd_data_out_0_246 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_246 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_247 <= 2'h0;
    end else if (bht_bank_sel_0_15_7) begin
      if (_T_8721) begin
        bht_bank_rd_data_out_0_247 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_247 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_248 <= 2'h0;
    end else if (bht_bank_sel_0_15_8) begin
      if (_T_8730) begin
        bht_bank_rd_data_out_0_248 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_248 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_249 <= 2'h0;
    end else if (bht_bank_sel_0_15_9) begin
      if (_T_8739) begin
        bht_bank_rd_data_out_0_249 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_249 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_250 <= 2'h0;
    end else if (bht_bank_sel_0_15_10) begin
      if (_T_8748) begin
        bht_bank_rd_data_out_0_250 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_250 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_251 <= 2'h0;
    end else if (bht_bank_sel_0_15_11) begin
      if (_T_8757) begin
        bht_bank_rd_data_out_0_251 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_251 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_252 <= 2'h0;
    end else if (bht_bank_sel_0_15_12) begin
      if (_T_8766) begin
        bht_bank_rd_data_out_0_252 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_252 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_253 <= 2'h0;
    end else if (bht_bank_sel_0_15_13) begin
      if (_T_8775) begin
        bht_bank_rd_data_out_0_253 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_253 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_254 <= 2'h0;
    end else if (bht_bank_sel_0_15_14) begin
      if (_T_8784) begin
        bht_bank_rd_data_out_0_254 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_254 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_255 <= 2'h0;
    end else if (bht_bank_sel_0_15_15) begin
      if (_T_8793) begin
        bht_bank_rd_data_out_0_255 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_255 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      exu_mp_way_f <= 1'h0;
    end else begin
      exu_mp_way_f <= io_exu_mp_pkt_way;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      exu_flush_final_d1 <= 1'h0;
    end else begin
      exu_flush_final_d1 <= io_exu_flush_final;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_lru_b0_f <= 256'h0;
    end else if (_T_213) begin
      btb_lru_b0_f <= btb_lru_b0_ns;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifc_fetch_adder_prior <= 31'h0;
    end else if (_T_373) begin
      ifc_fetch_adder_prior <= io_ifc_fetch_addr_f;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_0 <= 32'h0;
    end else if (rsenable_0) begin
      rets_out_0 <= rets_in_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_1 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_1 <= rets_in_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_2 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_2 <= rets_in_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_3 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_3 <= rets_in_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_4 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_4 <= rets_in_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_5 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_5 <= rets_in_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_6 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_6 <= rets_in_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_7 <= 32'h0;
    end else if (rs_push) begin
      rets_out_7 <= rets_out_6;
    end
  end
endmodule
