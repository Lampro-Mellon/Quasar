module sbox(
  input        clock,
  input        reset,
  input  [3:0] io_in,
  input        io_op,
  output       io_s_box_out_valid,
  output [3:0] io_s_box_out_bits,
  output       io_inv_s_box_out_valid,
  output [3:0] io_inv_s_box_out_bits
);
  wire  _T_1 = io_in == 4'h0; // @[quasar_wrapper.scala 185:74]
  wire  _T_3 = io_in == 4'h1; // @[quasar_wrapper.scala 185:74]
  wire  _T_5 = io_in == 4'h2; // @[quasar_wrapper.scala 185:74]
  wire  _T_7 = io_in == 4'h3; // @[quasar_wrapper.scala 185:74]
  wire  _T_9 = io_in == 4'h4; // @[quasar_wrapper.scala 185:74]
  wire  _T_11 = io_in == 4'h5; // @[quasar_wrapper.scala 185:74]
  wire  _T_13 = io_in == 4'h6; // @[quasar_wrapper.scala 185:74]
  wire  _T_15 = io_in == 4'h7; // @[quasar_wrapper.scala 185:74]
  wire  _T_17 = io_in == 4'h8; // @[quasar_wrapper.scala 185:74]
  wire  _T_19 = io_in == 4'h9; // @[quasar_wrapper.scala 185:74]
  wire  _T_21 = io_in == 4'ha; // @[quasar_wrapper.scala 185:74]
  wire  _T_23 = io_in == 4'hb; // @[quasar_wrapper.scala 185:74]
  wire  _T_25 = io_in == 4'hc; // @[quasar_wrapper.scala 185:74]
  wire  _T_27 = io_in == 4'hd; // @[quasar_wrapper.scala 185:74]
  wire  _T_29 = io_in == 4'he; // @[quasar_wrapper.scala 185:74]
  wire  _T_31 = io_in == 4'hf; // @[quasar_wrapper.scala 185:74]
  wire [2:0] _T_33 = _T_1 ? 3'h7 : 3'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_34 = _T_3 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_35 = _T_5 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_36 = _T_7 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_38 = _T_11 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_39 = _T_13 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_41 = _T_17 ? 3'h5 : 3'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_42 = _T_19 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_43 = _T_21 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_44 = _T_23 ? 3'h4 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_45 = _T_25 ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_46 = _T_27 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_47 = _T_29 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_48 = _T_31 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [2:0] _GEN_0 = {{1'd0}, _T_34}; // @[Mux.scala 27:72]
  wire [2:0] _T_49 = _T_33 | _GEN_0; // @[Mux.scala 27:72]
  wire [3:0] _GEN_1 = {{1'd0}, _T_49}; // @[Mux.scala 27:72]
  wire [3:0] _T_50 = _GEN_1 | _T_35; // @[Mux.scala 27:72]
  wire [3:0] _T_51 = _T_50 | _T_36; // @[Mux.scala 27:72]
  wire [3:0] _T_53 = _T_51 | _T_38; // @[Mux.scala 27:72]
  wire [3:0] _T_54 = _T_53 | _T_39; // @[Mux.scala 27:72]
  wire [3:0] _GEN_2 = {{3'd0}, _T_15}; // @[Mux.scala 27:72]
  wire [3:0] _T_55 = _T_54 | _GEN_2; // @[Mux.scala 27:72]
  wire [3:0] _GEN_3 = {{1'd0}, _T_41}; // @[Mux.scala 27:72]
  wire [3:0] _T_56 = _T_55 | _GEN_3; // @[Mux.scala 27:72]
  wire [3:0] _T_57 = _T_56 | _T_42; // @[Mux.scala 27:72]
  wire [3:0] _T_58 = _T_57 | _T_43; // @[Mux.scala 27:72]
  wire [3:0] _GEN_4 = {{1'd0}, _T_44}; // @[Mux.scala 27:72]
  wire [3:0] _T_59 = _T_58 | _GEN_4; // @[Mux.scala 27:72]
  wire [3:0] _GEN_5 = {{1'd0}, _T_45}; // @[Mux.scala 27:72]
  wire [3:0] _T_60 = _T_59 | _GEN_5; // @[Mux.scala 27:72]
  wire [3:0] _GEN_6 = {{2'd0}, _T_46}; // @[Mux.scala 27:72]
  wire [3:0] _T_61 = _T_60 | _GEN_6; // @[Mux.scala 27:72]
  wire [3:0] _T_62 = _T_61 | _T_47; // @[Mux.scala 27:72]
  wire [2:0] _T_97 = _T_1 ? 3'h4 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_98 = _T_3 ? 3'h7 : 3'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_99 = _T_5 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_101 = _T_9 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_102 = _T_11 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_103 = _T_13 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_105 = _T_17 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_106 = _T_19 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_107 = _T_21 ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_108 = _T_23 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_109 = _T_25 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_110 = _T_27 ? 3'h5 : 3'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_111 = _T_29 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_112 = _T_31 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_113 = _T_97 | _T_98; // @[Mux.scala 27:72]
  wire [3:0] _GEN_7 = {{1'd0}, _T_113}; // @[Mux.scala 27:72]
  wire [3:0] _T_114 = _GEN_7 | _T_99; // @[Mux.scala 27:72]
  wire [3:0] _GEN_8 = {{3'd0}, _T_7}; // @[Mux.scala 27:72]
  wire [3:0] _T_115 = _T_114 | _GEN_8; // @[Mux.scala 27:72]
  wire [3:0] _T_116 = _T_115 | _T_101; // @[Mux.scala 27:72]
  wire [3:0] _T_117 = _T_116 | _T_102; // @[Mux.scala 27:72]
  wire [3:0] _T_118 = _T_117 | _T_103; // @[Mux.scala 27:72]
  wire [3:0] _T_120 = _T_118 | _T_105; // @[Mux.scala 27:72]
  wire [3:0] _GEN_9 = {{2'd0}, _T_106}; // @[Mux.scala 27:72]
  wire [3:0] _T_121 = _T_120 | _GEN_9; // @[Mux.scala 27:72]
  wire [3:0] _GEN_10 = {{1'd0}, _T_107}; // @[Mux.scala 27:72]
  wire [3:0] _T_122 = _T_121 | _GEN_10; // @[Mux.scala 27:72]
  wire [3:0] _T_123 = _T_122 | _T_108; // @[Mux.scala 27:72]
  wire [3:0] _T_124 = _T_123 | _T_109; // @[Mux.scala 27:72]
  wire [3:0] _GEN_11 = {{1'd0}, _T_110}; // @[Mux.scala 27:72]
  wire [3:0] _T_125 = _T_124 | _GEN_11; // @[Mux.scala 27:72]
  wire [3:0] _GEN_12 = {{2'd0}, _T_111}; // @[Mux.scala 27:72]
  wire [3:0] _T_126 = _T_125 | _GEN_12; // @[Mux.scala 27:72]
  assign io_s_box_out_valid = ~io_op; // @[quasar_wrapper.scala 183:29]
  assign io_s_box_out_bits = _T_62 | _T_48; // @[quasar_wrapper.scala 185:21]
  assign io_inv_s_box_out_valid = io_op; // @[quasar_wrapper.scala 184:29]
  assign io_inv_s_box_out_bits = _T_126 | _T_112; // @[quasar_wrapper.scala 186:25]
endmodule
