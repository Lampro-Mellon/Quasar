module rvecc_encode_64(
  input  [63:0] io_din,
  output [6:0]  io_ecc_out
);
  wire  w0_0 = io_din[0]; // @[el2_lib.scala 343:39]
  wire  w0_1 = io_din[1]; // @[el2_lib.scala 343:39]
  wire  w1_1 = io_din[2]; // @[el2_lib.scala 344:39]
  wire  w0_2 = io_din[3]; // @[el2_lib.scala 343:39]
  wire  w0_3 = io_din[4]; // @[el2_lib.scala 343:39]
  wire  w1_3 = io_din[5]; // @[el2_lib.scala 344:39]
  wire  w0_4 = io_din[6]; // @[el2_lib.scala 343:39]
  wire  w2_3 = io_din[7]; // @[el2_lib.scala 345:39]
  wire  w0_5 = io_din[8]; // @[el2_lib.scala 343:39]
  wire  w1_5 = io_din[9]; // @[el2_lib.scala 344:39]
  wire  w0_6 = io_din[10]; // @[el2_lib.scala 343:39]
  wire  w0_7 = io_din[11]; // @[el2_lib.scala 343:39]
  wire  w1_7 = io_din[12]; // @[el2_lib.scala 344:39]
  wire  w0_8 = io_din[13]; // @[el2_lib.scala 343:39]
  wire  w2_7 = io_din[14]; // @[el2_lib.scala 345:39]
  wire  w0_9 = io_din[15]; // @[el2_lib.scala 343:39]
  wire  w1_9 = io_din[16]; // @[el2_lib.scala 344:39]
  wire  w0_10 = io_din[17]; // @[el2_lib.scala 343:39]
  wire  w3_7 = io_din[18]; // @[el2_lib.scala 346:39]
  wire  w0_11 = io_din[19]; // @[el2_lib.scala 343:39]
  wire  w1_11 = io_din[20]; // @[el2_lib.scala 344:39]
  wire  w0_12 = io_din[21]; // @[el2_lib.scala 343:39]
  wire  w2_11 = io_din[22]; // @[el2_lib.scala 345:39]
  wire  w0_13 = io_din[23]; // @[el2_lib.scala 343:39]
  wire  w1_13 = io_din[24]; // @[el2_lib.scala 344:39]
  wire  w0_14 = io_din[25]; // @[el2_lib.scala 343:39]
  wire  w0_15 = io_din[26]; // @[el2_lib.scala 343:39]
  wire  w1_15 = io_din[27]; // @[el2_lib.scala 344:39]
  wire  w0_16 = io_din[28]; // @[el2_lib.scala 343:39]
  wire  w2_15 = io_din[29]; // @[el2_lib.scala 345:39]
  wire  w0_17 = io_din[30]; // @[el2_lib.scala 343:39]
  wire  w1_17 = io_din[31]; // @[el2_lib.scala 344:39]
  wire  w0_18 = io_din[32]; // @[el2_lib.scala 343:39]
  wire  w3_15 = io_din[33]; // @[el2_lib.scala 346:39]
  wire  w0_19 = io_din[34]; // @[el2_lib.scala 343:39]
  wire  w1_19 = io_din[35]; // @[el2_lib.scala 344:39]
  wire  w0_20 = io_din[36]; // @[el2_lib.scala 343:39]
  wire  w2_19 = io_din[37]; // @[el2_lib.scala 345:39]
  wire  w0_21 = io_din[38]; // @[el2_lib.scala 343:39]
  wire  w1_21 = io_din[39]; // @[el2_lib.scala 344:39]
  wire  w0_22 = io_din[40]; // @[el2_lib.scala 343:39]
  wire  w4_15 = io_din[41]; // @[el2_lib.scala 347:39]
  wire  w0_23 = io_din[42]; // @[el2_lib.scala 343:39]
  wire  w1_23 = io_din[43]; // @[el2_lib.scala 344:39]
  wire  w0_24 = io_din[44]; // @[el2_lib.scala 343:39]
  wire  w2_23 = io_din[45]; // @[el2_lib.scala 345:39]
  wire  w0_25 = io_din[46]; // @[el2_lib.scala 343:39]
  wire  w1_25 = io_din[47]; // @[el2_lib.scala 344:39]
  wire  w0_26 = io_din[48]; // @[el2_lib.scala 343:39]
  wire  w3_23 = io_din[49]; // @[el2_lib.scala 346:39]
  wire  w0_27 = io_din[50]; // @[el2_lib.scala 343:39]
  wire  w1_27 = io_din[51]; // @[el2_lib.scala 344:39]
  wire  w0_28 = io_din[52]; // @[el2_lib.scala 343:39]
  wire  w2_27 = io_din[53]; // @[el2_lib.scala 345:39]
  wire  w0_29 = io_din[54]; // @[el2_lib.scala 343:39]
  wire  w1_29 = io_din[55]; // @[el2_lib.scala 344:39]
  wire  w0_30 = io_din[56]; // @[el2_lib.scala 343:39]
  wire  w0_31 = io_din[57]; // @[el2_lib.scala 343:39]
  wire  w1_31 = io_din[58]; // @[el2_lib.scala 344:39]
  wire  w0_32 = io_din[59]; // @[el2_lib.scala 343:39]
  wire  w2_31 = io_din[60]; // @[el2_lib.scala 345:39]
  wire  w0_33 = io_din[61]; // @[el2_lib.scala 343:39]
  wire  w1_33 = io_din[62]; // @[el2_lib.scala 344:39]
  wire  w0_34 = io_din[63]; // @[el2_lib.scala 343:39]
  wire [6:0] _T_210 = {w0_34,w1_33,w0_33,w2_31,w0_32,w1_31,w0_31}; // @[el2_lib.scala 351:27]
  wire  _T_211 = ^_T_210; // @[el2_lib.scala 351:34]
  wire [6:0] _T_217 = {w0_18,w1_17,w0_17,w2_15,w0_16,w1_15,w0_15}; // @[el2_lib.scala 351:44]
  wire [7:0] _T_224 = {w0_22,w1_21,w0_21,w2_19,w0_20,w1_19,w0_19,w3_15}; // @[el2_lib.scala 351:44]
  wire [14:0] _T_225 = {w0_22,w1_21,w0_21,w2_19,w0_20,w1_19,w0_19,w3_15,_T_217}; // @[el2_lib.scala 351:44]
  wire [7:0] _T_232 = {w0_26,w1_25,w0_25,w2_23,w0_24,w1_23,w0_23,w4_15}; // @[el2_lib.scala 351:44]
  wire [30:0] _T_241 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_232,_T_225}; // @[el2_lib.scala 351:44]
  wire  _T_242 = ^_T_241; // @[el2_lib.scala 351:51]
  wire [6:0] _T_248 = {w0_10,w1_9,w0_9,w2_7,w0_8,w1_7,w0_7}; // @[el2_lib.scala 351:61]
  wire [14:0] _T_256 = {w0_14,w1_13,w0_13,w2_11,w0_12,w1_11,w0_11,w3_7,_T_248}; // @[el2_lib.scala 351:61]
  wire [30:0] _T_272 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_232,_T_256}; // @[el2_lib.scala 351:61]
  wire  _T_273 = ^_T_272; // @[el2_lib.scala 351:68]
  wire [6:0] _T_279 = {w0_6,w1_5,w0_5,w2_3,w0_4,w1_3,w0_3}; // @[el2_lib.scala 351:78]
  wire [14:0] _T_287 = {w0_14,w1_13,w0_13,w2_11,w0_12,w1_11,w0_11,w3_7,_T_279}; // @[el2_lib.scala 351:78]
  wire [30:0] _T_303 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_224,_T_287}; // @[el2_lib.scala 351:78]
  wire  _T_304 = ^_T_303; // @[el2_lib.scala 351:85]
  wire [7:0] _T_311 = {w2_7,w0_6,w1_5,w0_5,w2_3,w0_2,w1_1,w0_1}; // @[el2_lib.scala 351:95]
  wire [16:0] _T_320 = {w0_17,w2_15,w0_14,w1_13,w0_13,w2_11,w0_10,w1_9,w0_9,_T_311}; // @[el2_lib.scala 351:95]
  wire [8:0] _T_328 = {w1_25,w0_25,w2_23,w0_22,w1_21,w0_21,w2_19,w0_18,w1_17}; // @[el2_lib.scala 351:95]
  wire [17:0] _T_337 = {w0_34,w1_33,w0_33,w2_31,w0_30,w1_29,w0_29,w2_27,w0_26,_T_328}; // @[el2_lib.scala 351:95]
  wire [34:0] _T_338 = {_T_337,_T_320}; // @[el2_lib.scala 351:95]
  wire  _T_339 = ^_T_338; // @[el2_lib.scala 351:102]
  wire [7:0] _T_346 = {w1_7,w0_6,w1_5,w0_4,w1_3,w0_2,w1_1,w0_0}; // @[el2_lib.scala 351:112]
  wire [16:0] _T_355 = {w0_16,w1_15,w0_14,w1_13,w0_12,w1_11,w0_10,w1_9,w0_8,_T_346}; // @[el2_lib.scala 351:112]
  wire [8:0] _T_363 = {w1_25,w0_24,w1_23,w0_22,w1_21,w0_20,w1_19,w0_18,w1_17}; // @[el2_lib.scala 351:112]
  wire [17:0] _T_372 = {w0_34,w1_33,w0_32,w1_31,w0_30,w1_29,w0_28,w1_27,w0_26,_T_363}; // @[el2_lib.scala 351:112]
  wire [34:0] _T_373 = {_T_372,_T_355}; // @[el2_lib.scala 351:112]
  wire  _T_374 = ^_T_373; // @[el2_lib.scala 351:119]
  wire [7:0] _T_381 = {w0_7,w0_6,w0_5,w0_4,w0_3,w0_2,w0_1,w0_0}; // @[el2_lib.scala 351:129]
  wire [16:0] _T_390 = {w0_16,w0_15,w0_14,w0_13,w0_12,w0_11,w0_10,w0_9,w0_8,_T_381}; // @[el2_lib.scala 351:129]
  wire [8:0] _T_398 = {w0_25,w0_24,w0_23,w0_22,w0_21,w0_20,w0_19,w0_18,w0_17}; // @[el2_lib.scala 351:129]
  wire [17:0] _T_407 = {w0_34,w0_33,w0_32,w0_31,w0_30,w0_29,w0_28,w0_27,w0_26,_T_398}; // @[el2_lib.scala 351:129]
  wire [34:0] _T_408 = {_T_407,_T_390}; // @[el2_lib.scala 351:129]
  wire  _T_409 = ^_T_408; // @[el2_lib.scala 351:136]
  wire [2:0] _T_411 = {_T_339,_T_374,_T_409}; // @[Cat.scala 29:58]
  wire [3:0] _T_414 = {_T_211,_T_242,_T_273,_T_304}; // @[Cat.scala 29:58]
  assign io_ecc_out = {_T_414,_T_411}; // @[el2_lib.scala 351:16]
endmodule
module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [95:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [63:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] m1_io_din; // @[el2_ifu_mem_ctl.scala 342:18]
  wire [6:0] m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 342:18]
  wire [63:0] m2_io_din; // @[el2_ifu_mem_ctl.scala 343:18]
  wire [6:0] m2_io_ecc_out; // @[el2_ifu_mem_ctl.scala 343:18]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 184:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 320:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 321:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 321:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 253:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 553:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 555:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 186:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 308:34]
  wire [4:0] _GEN_464 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 670:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_464 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 670:53]
  wire [1:0] _GEN_465 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 673:91]
  wire [1:0] _T_2277 = ic_fetch_val_shift_right[3:2] & _GEN_465; // @[el2_ifu_mem_ctl.scala 673:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 322:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 275:46]
  wire [1:0] _GEN_466 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 673:113]
  wire [1:0] _T_2278 = _T_2277 & _GEN_466; // @[el2_ifu_mem_ctl.scala 673:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 659:59]
  wire [1:0] _GEN_467 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 673:130]
  wire [1:0] _T_2279 = _T_2278 | _GEN_467; // @[el2_ifu_mem_ctl.scala 673:130]
  wire  _T_2280 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 673:154]
  wire [1:0] _GEN_468 = {{1'd0}, _T_2280}; // @[el2_ifu_mem_ctl.scala 673:152]
  wire [1:0] _T_2281 = _T_2279 & _GEN_468; // @[el2_ifu_mem_ctl.scala 673:152]
  wire [1:0] _T_2270 = ic_fetch_val_shift_right[1:0] & _GEN_465; // @[el2_ifu_mem_ctl.scala 673:91]
  wire [1:0] _T_2271 = _T_2270 & _GEN_466; // @[el2_ifu_mem_ctl.scala 673:113]
  wire [1:0] _T_2272 = _T_2271 | _GEN_467; // @[el2_ifu_mem_ctl.scala 673:130]
  wire [1:0] _T_2274 = _T_2272 & _GEN_468; // @[el2_ifu_mem_ctl.scala 673:152]
  wire [3:0] iccm_ecc_word_enable = {_T_2281,_T_2274}; // @[Cat.scala 29:58]
  wire  _T_2381 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_2382 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_2383 = _T_2381 ^ _T_2382; // @[el2_lib.scala 301:35]
  wire [5:0] _T_2391 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_2392 = ^_T_2391; // @[el2_lib.scala 301:83]
  wire  _T_2393 = io_iccm_rd_data_ecc[37] ^ _T_2392; // @[el2_lib.scala 301:71]
  wire [6:0] _T_2400 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_2408 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_2400}; // @[el2_lib.scala 301:103]
  wire  _T_2409 = ^_T_2408; // @[el2_lib.scala 301:110]
  wire  _T_2410 = io_iccm_rd_data_ecc[36] ^ _T_2409; // @[el2_lib.scala 301:98]
  wire [6:0] _T_2417 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_2425 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_2417}; // @[el2_lib.scala 301:130]
  wire  _T_2426 = ^_T_2425; // @[el2_lib.scala 301:137]
  wire  _T_2427 = io_iccm_rd_data_ecc[35] ^ _T_2426; // @[el2_lib.scala 301:125]
  wire [8:0] _T_2436 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_2445 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_2436}; // @[el2_lib.scala 301:157]
  wire  _T_2446 = ^_T_2445; // @[el2_lib.scala 301:164]
  wire  _T_2447 = io_iccm_rd_data_ecc[34] ^ _T_2446; // @[el2_lib.scala 301:152]
  wire [8:0] _T_2456 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_2465 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_2456}; // @[el2_lib.scala 301:184]
  wire  _T_2466 = ^_T_2465; // @[el2_lib.scala 301:191]
  wire  _T_2467 = io_iccm_rd_data_ecc[33] ^ _T_2466; // @[el2_lib.scala 301:179]
  wire [8:0] _T_2476 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_2485 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_2476}; // @[el2_lib.scala 301:211]
  wire  _T_2486 = ^_T_2485; // @[el2_lib.scala 301:218]
  wire  _T_2487 = io_iccm_rd_data_ecc[32] ^ _T_2486; // @[el2_lib.scala 301:206]
  wire [6:0] _T_2493 = {_T_2383,_T_2393,_T_2410,_T_2427,_T_2447,_T_2467,_T_2487}; // @[Cat.scala 29:58]
  wire  _T_2494 = _T_2493 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_2495 = iccm_ecc_word_enable[0] & _T_2494; // @[el2_lib.scala 302:32]
  wire  _T_2497 = _T_2495 & _T_2493[6]; // @[el2_lib.scala 302:53]
  wire  _T_2766 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_2767 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_2768 = _T_2766 ^ _T_2767; // @[el2_lib.scala 301:35]
  wire [5:0] _T_2776 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_2777 = ^_T_2776; // @[el2_lib.scala 301:83]
  wire  _T_2778 = io_iccm_rd_data_ecc[76] ^ _T_2777; // @[el2_lib.scala 301:71]
  wire [6:0] _T_2785 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_2793 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_2785}; // @[el2_lib.scala 301:103]
  wire  _T_2794 = ^_T_2793; // @[el2_lib.scala 301:110]
  wire  _T_2795 = io_iccm_rd_data_ecc[75] ^ _T_2794; // @[el2_lib.scala 301:98]
  wire [6:0] _T_2802 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_2810 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_2802}; // @[el2_lib.scala 301:130]
  wire  _T_2811 = ^_T_2810; // @[el2_lib.scala 301:137]
  wire  _T_2812 = io_iccm_rd_data_ecc[74] ^ _T_2811; // @[el2_lib.scala 301:125]
  wire [8:0] _T_2821 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_2830 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_2821}; // @[el2_lib.scala 301:157]
  wire  _T_2831 = ^_T_2830; // @[el2_lib.scala 301:164]
  wire  _T_2832 = io_iccm_rd_data_ecc[73] ^ _T_2831; // @[el2_lib.scala 301:152]
  wire [8:0] _T_2841 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_2850 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_2841}; // @[el2_lib.scala 301:184]
  wire  _T_2851 = ^_T_2850; // @[el2_lib.scala 301:191]
  wire  _T_2852 = io_iccm_rd_data_ecc[72] ^ _T_2851; // @[el2_lib.scala 301:179]
  wire [8:0] _T_2861 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_2870 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_2861}; // @[el2_lib.scala 301:211]
  wire  _T_2871 = ^_T_2870; // @[el2_lib.scala 301:218]
  wire  _T_2872 = io_iccm_rd_data_ecc[71] ^ _T_2871; // @[el2_lib.scala 301:206]
  wire [6:0] _T_2878 = {_T_2768,_T_2778,_T_2795,_T_2812,_T_2832,_T_2852,_T_2872}; // @[Cat.scala 29:58]
  wire  _T_2879 = _T_2878 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_2880 = iccm_ecc_word_enable[1] & _T_2879; // @[el2_lib.scala 302:32]
  wire  _T_2882 = _T_2880 & _T_2878[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_2497,_T_2882}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 189:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 637:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 190:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 191:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 482:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 191:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 191:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 191:72]
  wire  _T_1646 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1651 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1671 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 532:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 396:42]
  wire  _T_1673 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 532:79]
  wire  _T_1674 = _T_1671 | _T_1673; // @[el2_ifu_mem_ctl.scala 532:56]
  wire  _T_1675 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 532:122]
  wire  _T_1676 = ~_T_1675; // @[el2_ifu_mem_ctl.scala 532:101]
  wire  _T_1677 = _T_1674 & _T_1676; // @[el2_ifu_mem_ctl.scala 532:99]
  wire  _T_1678 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1692 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 539:45]
  wire  _T_1693 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 539:69]
  wire  _T_1694 = _T_1692 & _T_1693; // @[el2_ifu_mem_ctl.scala 539:67]
  wire  _T_1695 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_55 = _T_1678 ? _T_1694 : _T_1695; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_1651 ? _T_1677 : _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_1646 ? 1'h0 : _GEN_59; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 191:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 193:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 193:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 283:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 283:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 705:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 283:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 274:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 274:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 324:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 274:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 274:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 283:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 283:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 283:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 283:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 552:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 594:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 621:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 310:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 602:56]
  wire  _T_1797 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 619:69]
  wire  _T_1798 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 619:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_1797 : _T_1798; // @[el2_ifu_mem_ctl.scala 619:28]
  wire  _T_1744 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 598:68]
  wire  _T_1745 = ic_act_miss_f | _T_1744; // @[el2_ifu_mem_ctl.scala 598:48]
  wire  bus_reset_data_beat_cnt = _T_1745 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 598:91]
  wire  _T_1741 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 597:50]
  wire  _T_1742 = bus_ifu_wr_en_ff & _T_1741; // @[el2_ifu_mem_ctl.scala 597:48]
  wire  _T_1743 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 597:72]
  wire  bus_inc_data_beat_cnt = _T_1742 & _T_1743; // @[el2_ifu_mem_ctl.scala 597:70]
  wire [2:0] _T_1749 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 601:115]
  wire [2:0] _T_1751 = bus_inc_data_beat_cnt ? _T_1749 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_1746 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 599:32]
  wire  _T_1747 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 599:57]
  wire  bus_hold_data_beat_cnt = _T_1746 & _T_1747; // @[el2_ifu_mem_ctl.scala 599:55]
  wire [2:0] _T_1752 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_1751 | _T_1752; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 193:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 193:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 194:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 193:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 194:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 200:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 200:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 432:45]
  wire  _T_1276 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 453:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 409:60]
  wire  _T_1307 = _T_1276 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1280 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 453:127]
  wire  _T_1308 = _T_1280 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1315 = _T_1307 | _T_1308; // @[Mux.scala 27:72]
  wire  _T_1284 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 453:127]
  wire  _T_1309 = _T_1284 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1316 = _T_1315 | _T_1309; // @[Mux.scala 27:72]
  wire  _T_1288 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 453:127]
  wire  _T_1310 = _T_1288 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1317 = _T_1316 | _T_1310; // @[Mux.scala 27:72]
  wire  _T_1292 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 453:127]
  wire  _T_1311 = _T_1292 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1318 = _T_1317 | _T_1311; // @[Mux.scala 27:72]
  wire  _T_1296 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 453:127]
  wire  _T_1312 = _T_1296 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1319 = _T_1318 | _T_1312; // @[Mux.scala 27:72]
  wire  _T_1300 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 453:127]
  wire  _T_1313 = _T_1300 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1320 = _T_1319 | _T_1313; // @[Mux.scala 27:72]
  wire  _T_1304 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 453:127]
  wire  _T_1314 = _T_1304 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_1320 | _T_1314; // @[Mux.scala 27:72]
  wire  _T_1362 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 455:69]
  wire  _T_1363 = ic_miss_buff_data_valid_bypass_index & _T_1362; // @[el2_ifu_mem_ctl.scala 455:67]
  wire  _T_1365 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 455:91]
  wire  _T_1366 = _T_1363 & _T_1365; // @[el2_ifu_mem_ctl.scala 455:89]
  wire  _T_1371 = _T_1363 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 456:65]
  wire  _T_1372 = _T_1366 | _T_1371; // @[el2_ifu_mem_ctl.scala 455:112]
  wire  _T_1374 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 457:43]
  wire  _T_1377 = _T_1374 & _T_1365; // @[el2_ifu_mem_ctl.scala 457:65]
  wire  _T_1378 = _T_1372 | _T_1377; // @[el2_ifu_mem_ctl.scala 456:88]
  wire  _T_1382 = _T_1374 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 458:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 435:75]
  wire  _T_1322 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 454:110]
  wire  _T_1346 = _T_1322 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1325 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 454:110]
  wire  _T_1347 = _T_1325 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1354 = _T_1346 | _T_1347; // @[Mux.scala 27:72]
  wire  _T_1328 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 454:110]
  wire  _T_1348 = _T_1328 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1355 = _T_1354 | _T_1348; // @[Mux.scala 27:72]
  wire  _T_1331 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 454:110]
  wire  _T_1349 = _T_1331 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1356 = _T_1355 | _T_1349; // @[Mux.scala 27:72]
  wire  _T_1334 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 454:110]
  wire  _T_1350 = _T_1334 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1357 = _T_1356 | _T_1350; // @[Mux.scala 27:72]
  wire  _T_1337 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 454:110]
  wire  _T_1351 = _T_1337 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1358 = _T_1357 | _T_1351; // @[Mux.scala 27:72]
  wire  _T_1340 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 454:110]
  wire  _T_1352 = _T_1340 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1359 = _T_1358 | _T_1352; // @[Mux.scala 27:72]
  wire  _T_1343 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 454:110]
  wire  _T_1353 = _T_1343 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_1359 | _T_1353; // @[Mux.scala 27:72]
  wire  _T_1383 = _T_1382 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 458:87]
  wire  _T_1384 = _T_1378 | _T_1383; // @[el2_ifu_mem_ctl.scala 457:88]
  wire  _T_1388 = ic_miss_buff_data_valid_bypass_index & _T_1304; // @[el2_ifu_mem_ctl.scala 459:43]
  wire  miss_buff_hit_unq_f = _T_1384 | _T_1388; // @[el2_ifu_mem_ctl.scala 458:131]
  wire  _T_1404 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 464:55]
  wire  _T_1405 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 464:87]
  wire  _T_1406 = _T_1404 | _T_1405; // @[el2_ifu_mem_ctl.scala 464:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_1406; // @[el2_ifu_mem_ctl.scala 464:41]
  wire  _T_1389 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 461:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 311:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[6]; // @[el2_ifu_mem_ctl.scala 452:51]
  wire  _T_1390 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 461:68]
  wire  _T_1391 = miss_buff_hit_unq_f & _T_1390; // @[el2_ifu_mem_ctl.scala 461:66]
  wire  stream_hit_f = _T_1389 & _T_1391; // @[el2_ifu_mem_ctl.scala 461:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 278:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 278:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 278:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 604:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 631:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 204:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 204:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 204:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 204:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 204:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 205:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 205:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 205:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 206:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 206:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 206:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 207:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 208:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 208:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 208:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 196:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 208:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 208:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 208:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 209:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 209:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 209:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 209:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 210:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 211:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 211:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 211:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 210:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 209:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 208:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 207:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 206:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 205:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 204:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_1401 = byp_fetch_index[4:1] == 4'h7; // @[el2_ifu_mem_ctl.scala 463:60]
  wire  _T_1402 = _T_1401 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 463:92]
  wire  stream_eol_f = _T_1402 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 463:110]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 219:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 219:87]
  wire  _T_113 = _T_111 & _T_1743; // @[el2_ifu_mem_ctl.scala 219:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 219:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 223:48]
  wire  _T_126 = _T_124 & _T_1743; // @[el2_ifu_mem_ctl.scala 223:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 223:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 284:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 284:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 284:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 284:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 285:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 284:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 285:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 338:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 285:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 285:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 285:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 227:50]
  wire  _T_137 = _T_135 & _T_1743; // @[el2_ifu_mem_ctl.scala 227:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 286:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 287:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 287:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 286:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 228:35]
  wire  _T_143 = _T_141 & _T_1743; // @[el2_ifu_mem_ctl.scala 228:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 228:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 227:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 233:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 232:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 232:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 237:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 237:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 194:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 194:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 194:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 194:91]
  wire  _T_30 = ic_act_miss_f & _T_1743; // @[el2_ifu_mem_ctl.scala 201:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 212:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 212:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 212:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 212:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 212:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 212:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 216:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 216:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 216:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 220:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 220:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 224:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 224:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 229:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 229:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 229:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 234:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 234:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 254:95]
  wire  _T_175 = _T_1404 & _T_174; // @[el2_ifu_mem_ctl.scala 254:93]
  wire  crit_wd_byp_ok_ff = _T_1405 | _T_175; // @[el2_ifu_mem_ctl.scala 254:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 255:36]
  wire  _T_180 = _T_1404 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 255:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 255:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 255:70]
  wire  _T_184 = _T_1404 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 256:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 256:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 255:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 256:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 257:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 257:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 256:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 259:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 259:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:35]
  reg [6:0] _T_4322; // @[el2_ifu_mem_ctl.scala 733:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_4322[5:0]; // @[el2_ifu_mem_ctl.scala 732:27]
  wire [6:0] _GEN_473 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 729:121]
  wire  _T_4187 = _GEN_473 == 7'h7f; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4189 = _T_4187 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3678; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_3678[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_474 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4190 = _T_4189 & _GEN_474; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4183 = _GEN_473 == 7'h7e; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4185 = _T_4183 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3674; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_3674[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_476 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4186 = _T_4185 & _GEN_476; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4179 = _GEN_473 == 7'h7d; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4181 = _T_4179 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3670; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_3670[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_478 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4182 = _T_4181 & _GEN_478; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4175 = _GEN_473 == 7'h7c; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4177 = _T_4175 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3666; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_3666[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_480 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4178 = _T_4177 & _GEN_480; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4171 = _GEN_473 == 7'h7b; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4173 = _T_4171 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3662; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_3662[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_482 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4174 = _T_4173 & _GEN_482; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4167 = _GEN_473 == 7'h7a; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4169 = _T_4167 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3658; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_3658[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_484 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4170 = _T_4169 & _GEN_484; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4163 = _GEN_473 == 7'h79; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4165 = _T_4163 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3654; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_3654[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_486 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4166 = _T_4165 & _GEN_486; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4159 = _GEN_473 == 7'h78; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4161 = _T_4159 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3650; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_3650[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_488 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4162 = _T_4161 & _GEN_488; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4155 = _GEN_473 == 7'h77; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4157 = _T_4155 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3646; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_3646[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_490 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4158 = _T_4157 & _GEN_490; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4151 = _GEN_473 == 7'h76; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4153 = _T_4151 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3642; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_3642[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_492 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4154 = _T_4153 & _GEN_492; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [59:0] _T_4199 = {_T_4190,_T_4186,_T_4182,_T_4178,_T_4174,_T_4170,_T_4166,_T_4162,_T_4158,_T_4154}; // @[Cat.scala 29:58]
  wire  _T_4147 = _GEN_473 == 7'h75; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4149 = _T_4147 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3638; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_3638[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_494 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4150 = _T_4149 & _GEN_494; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4143 = _GEN_473 == 7'h74; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4145 = _T_4143 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3634; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_3634[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_496 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4146 = _T_4145 & _GEN_496; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4139 = _GEN_473 == 7'h73; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4141 = _T_4139 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3630; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_3630[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_498 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4142 = _T_4141 & _GEN_498; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4135 = _GEN_473 == 7'h72; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4137 = _T_4135 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3626; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_3626[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_500 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4138 = _T_4137 & _GEN_500; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4131 = _GEN_473 == 7'h71; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4133 = _T_4131 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3622; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_3622[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_502 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4134 = _T_4133 & _GEN_502; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4127 = _GEN_473 == 7'h70; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4129 = _T_4127 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3618; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_3618[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_504 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4130 = _T_4129 & _GEN_504; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4123 = _GEN_473 == 7'h6f; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4125 = _T_4123 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3614; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_3614[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_506 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4126 = _T_4125 & _GEN_506; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4119 = _GEN_473 == 7'h6e; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4121 = _T_4119 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3610; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_3610[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_508 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4122 = _T_4121 & _GEN_508; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4115 = _GEN_473 == 7'h6d; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4117 = _T_4115 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3606; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_3606[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_510 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4118 = _T_4117 & _GEN_510; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [113:0] _T_4208 = {_T_4199,_T_4150,_T_4146,_T_4142,_T_4138,_T_4134,_T_4130,_T_4126,_T_4122,_T_4118}; // @[Cat.scala 29:58]
  wire  _T_4111 = _GEN_473 == 7'h6c; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4113 = _T_4111 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3602; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_3602[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_512 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4114 = _T_4113 & _GEN_512; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4107 = _GEN_473 == 7'h6b; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4109 = _T_4107 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3598; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_3598[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_514 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4110 = _T_4109 & _GEN_514; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4103 = _GEN_473 == 7'h6a; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4105 = _T_4103 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3594; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_3594[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_516 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4106 = _T_4105 & _GEN_516; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4099 = _GEN_473 == 7'h69; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4101 = _T_4099 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3590; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_3590[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_518 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4102 = _T_4101 & _GEN_518; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4095 = _GEN_473 == 7'h68; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4097 = _T_4095 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3586; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_3586[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_520 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4098 = _T_4097 & _GEN_520; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4091 = _GEN_473 == 7'h67; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4093 = _T_4091 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3582; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_3582[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_522 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4094 = _T_4093 & _GEN_522; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4087 = _GEN_473 == 7'h66; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4089 = _T_4087 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3578; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_3578[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_524 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4090 = _T_4089 & _GEN_524; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4083 = _GEN_473 == 7'h65; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4085 = _T_4083 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3574; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_3574[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_526 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4086 = _T_4085 & _GEN_526; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4079 = _GEN_473 == 7'h64; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4081 = _T_4079 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3570; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_3570[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_528 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4082 = _T_4081 & _GEN_528; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [167:0] _T_4217 = {_T_4208,_T_4114,_T_4110,_T_4106,_T_4102,_T_4098,_T_4094,_T_4090,_T_4086,_T_4082}; // @[Cat.scala 29:58]
  wire  _T_4075 = _GEN_473 == 7'h63; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4077 = _T_4075 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3566; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_3566[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_530 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4078 = _T_4077 & _GEN_530; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4071 = _GEN_473 == 7'h62; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4073 = _T_4071 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3562; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_3562[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_532 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4074 = _T_4073 & _GEN_532; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4067 = _GEN_473 == 7'h61; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4069 = _T_4067 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3558; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_3558[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_534 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4070 = _T_4069 & _GEN_534; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4063 = _GEN_473 == 7'h60; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4065 = _T_4063 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3554; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_3554[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_536 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4066 = _T_4065 & _GEN_536; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4059 = _GEN_473 == 7'h5f; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4061 = _T_4059 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3550; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_3550[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_538 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4062 = _T_4061 & _GEN_538; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4055 = _GEN_473 == 7'h5e; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4057 = _T_4055 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3546; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_3546[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_540 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4058 = _T_4057 & _GEN_540; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4051 = _GEN_473 == 7'h5d; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4053 = _T_4051 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3542; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_3542[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_542 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4054 = _T_4053 & _GEN_542; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4047 = _GEN_473 == 7'h5c; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4049 = _T_4047 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3538; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_3538[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_544 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4050 = _T_4049 & _GEN_544; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4043 = _GEN_473 == 7'h5b; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4045 = _T_4043 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3534; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_3534[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_546 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4046 = _T_4045 & _GEN_546; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [221:0] _T_4226 = {_T_4217,_T_4078,_T_4074,_T_4070,_T_4066,_T_4062,_T_4058,_T_4054,_T_4050,_T_4046}; // @[Cat.scala 29:58]
  wire  _T_4039 = _GEN_473 == 7'h5a; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4041 = _T_4039 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3530; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_3530[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_548 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4042 = _T_4041 & _GEN_548; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4035 = _GEN_473 == 7'h59; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4037 = _T_4035 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3526; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_3526[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_550 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4038 = _T_4037 & _GEN_550; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4031 = _GEN_473 == 7'h58; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4033 = _T_4031 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3522; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_3522[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_552 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4034 = _T_4033 & _GEN_552; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4027 = _GEN_473 == 7'h57; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4029 = _T_4027 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3518; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_3518[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_554 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4030 = _T_4029 & _GEN_554; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4023 = _GEN_473 == 7'h56; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4025 = _T_4023 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3514; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_3514[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_556 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4026 = _T_4025 & _GEN_556; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4019 = _GEN_473 == 7'h55; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4021 = _T_4019 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3510; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_3510[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_558 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4022 = _T_4021 & _GEN_558; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4015 = _GEN_473 == 7'h54; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4017 = _T_4015 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3506; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_3506[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_560 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4018 = _T_4017 & _GEN_560; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4011 = _GEN_473 == 7'h53; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4013 = _T_4011 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3502; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_3502[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_562 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4014 = _T_4013 & _GEN_562; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_4007 = _GEN_473 == 7'h52; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4009 = _T_4007 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3498; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_3498[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_564 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4010 = _T_4009 & _GEN_564; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [275:0] _T_4235 = {_T_4226,_T_4042,_T_4038,_T_4034,_T_4030,_T_4026,_T_4022,_T_4018,_T_4014,_T_4010}; // @[Cat.scala 29:58]
  wire  _T_4003 = _GEN_473 == 7'h51; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4005 = _T_4003 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3494; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_3494[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_566 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4006 = _T_4005 & _GEN_566; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3999 = _GEN_473 == 7'h50; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_4001 = _T_3999 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3490; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_3490[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_568 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_4002 = _T_4001 & _GEN_568; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3995 = _GEN_473 == 7'h4f; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3997 = _T_3995 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3486; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_3486[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_570 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3998 = _T_3997 & _GEN_570; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3991 = _GEN_473 == 7'h4e; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3993 = _T_3991 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3482; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_3482[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_572 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3994 = _T_3993 & _GEN_572; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3987 = _GEN_473 == 7'h4d; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3989 = _T_3987 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3478; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_3478[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_574 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3990 = _T_3989 & _GEN_574; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3983 = _GEN_473 == 7'h4c; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3985 = _T_3983 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3474; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_3474[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_576 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3986 = _T_3985 & _GEN_576; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3979 = _GEN_473 == 7'h4b; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3981 = _T_3979 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3470; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_3470[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_578 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3982 = _T_3981 & _GEN_578; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3975 = _GEN_473 == 7'h4a; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3977 = _T_3975 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3466; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_3466[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_580 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3978 = _T_3977 & _GEN_580; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3971 = _GEN_473 == 7'h49; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3973 = _T_3971 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3462; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_3462[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_582 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3974 = _T_3973 & _GEN_582; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [329:0] _T_4244 = {_T_4235,_T_4006,_T_4002,_T_3998,_T_3994,_T_3990,_T_3986,_T_3982,_T_3978,_T_3974}; // @[Cat.scala 29:58]
  wire  _T_3967 = _GEN_473 == 7'h48; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3969 = _T_3967 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3458; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_3458[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_584 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3970 = _T_3969 & _GEN_584; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3963 = _GEN_473 == 7'h47; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3965 = _T_3963 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3454; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_3454[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_586 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3966 = _T_3965 & _GEN_586; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3959 = _GEN_473 == 7'h46; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3961 = _T_3959 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3450; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_3450[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_588 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3962 = _T_3961 & _GEN_588; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3955 = _GEN_473 == 7'h45; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3957 = _T_3955 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3446; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_3446[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_590 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3958 = _T_3957 & _GEN_590; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3951 = _GEN_473 == 7'h44; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3953 = _T_3951 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3442; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_3442[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_592 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3954 = _T_3953 & _GEN_592; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3947 = _GEN_473 == 7'h43; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3949 = _T_3947 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3438; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_3438[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_594 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3950 = _T_3949 & _GEN_594; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3943 = _GEN_473 == 7'h42; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3945 = _T_3943 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3434; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_3434[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_596 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3946 = _T_3945 & _GEN_596; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3939 = _GEN_473 == 7'h41; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3941 = _T_3939 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3430; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_3430[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_598 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3942 = _T_3941 & _GEN_598; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3935 = _GEN_473 == 7'h40; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3937 = _T_3935 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3426; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_3426[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3938 = _T_3937 & _GEN_600; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [383:0] _T_4253 = {_T_4244,_T_3970,_T_3966,_T_3962,_T_3958,_T_3954,_T_3950,_T_3946,_T_3942,_T_3938}; // @[Cat.scala 29:58]
  wire  _T_3931 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3933 = _T_3931 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3422; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_3422[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3934 = _T_3933 & _GEN_601; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3927 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3929 = _T_3927 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3418; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_3418[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3930 = _T_3929 & _GEN_602; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3923 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3925 = _T_3923 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3414; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_3414[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3926 = _T_3925 & _GEN_603; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3919 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3921 = _T_3919 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3410; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_3410[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3922 = _T_3921 & _GEN_604; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3915 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3917 = _T_3915 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3406; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_3406[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3918 = _T_3917 & _GEN_605; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3911 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3913 = _T_3911 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3402; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_3402[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3914 = _T_3913 & _GEN_606; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3907 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3909 = _T_3907 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3398; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_3398[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3910 = _T_3909 & _GEN_607; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3903 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3905 = _T_3903 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3394; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_3394[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3906 = _T_3905 & _GEN_608; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3899 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3901 = _T_3899 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3390; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_3390[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3902 = _T_3901 & _GEN_609; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [437:0] _T_4262 = {_T_4253,_T_3934,_T_3930,_T_3926,_T_3922,_T_3918,_T_3914,_T_3910,_T_3906,_T_3902}; // @[Cat.scala 29:58]
  wire  _T_3895 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3897 = _T_3895 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3386; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_3386[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3898 = _T_3897 & _GEN_610; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3891 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3893 = _T_3891 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3382; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_3382[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3894 = _T_3893 & _GEN_611; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3887 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3889 = _T_3887 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3378; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_3378[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3890 = _T_3889 & _GEN_612; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3883 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3885 = _T_3883 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3374; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_3374[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3886 = _T_3885 & _GEN_613; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3879 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3881 = _T_3879 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3370; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_3370[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3882 = _T_3881 & _GEN_614; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3875 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3877 = _T_3875 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3366; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_3366[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3878 = _T_3877 & _GEN_615; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3871 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3873 = _T_3871 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3362; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_3362[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3874 = _T_3873 & _GEN_616; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3867 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3869 = _T_3867 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3358; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_3358[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3870 = _T_3869 & _GEN_617; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3863 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3865 = _T_3863 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3354; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_3354[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3866 = _T_3865 & _GEN_618; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [491:0] _T_4271 = {_T_4262,_T_3898,_T_3894,_T_3890,_T_3886,_T_3882,_T_3878,_T_3874,_T_3870,_T_3866}; // @[Cat.scala 29:58]
  wire  _T_3859 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3861 = _T_3859 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3350; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_3350[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3862 = _T_3861 & _GEN_619; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3855 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3857 = _T_3855 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3346; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_3346[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3858 = _T_3857 & _GEN_620; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3851 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3853 = _T_3851 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3342; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_3342[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3854 = _T_3853 & _GEN_621; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3847 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3849 = _T_3847 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3338; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_3338[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3850 = _T_3849 & _GEN_622; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3843 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3845 = _T_3843 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3334; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_3334[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3846 = _T_3845 & _GEN_623; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3839 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3841 = _T_3839 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3330; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_3330[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3842 = _T_3841 & _GEN_624; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3835 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3837 = _T_3835 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3326; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_3326[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3838 = _T_3837 & _GEN_625; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3831 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3833 = _T_3831 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3322; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_3322[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3834 = _T_3833 & _GEN_626; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3827 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3829 = _T_3827 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3318; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_3318[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3830 = _T_3829 & _GEN_627; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [545:0] _T_4280 = {_T_4271,_T_3862,_T_3858,_T_3854,_T_3850,_T_3846,_T_3842,_T_3838,_T_3834,_T_3830}; // @[Cat.scala 29:58]
  wire  _T_3823 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3825 = _T_3823 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3314; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_3314[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3826 = _T_3825 & _GEN_628; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3819 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3821 = _T_3819 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3310; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_3310[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3822 = _T_3821 & _GEN_629; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3815 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3817 = _T_3815 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3306; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_3306[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3818 = _T_3817 & _GEN_630; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3811 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3813 = _T_3811 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3302; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_3302[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3814 = _T_3813 & _GEN_631; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3807 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3809 = _T_3807 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3298; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_3298[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3810 = _T_3809 & _GEN_632; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3803 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3805 = _T_3803 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3294; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_3294[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3806 = _T_3805 & _GEN_633; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3799 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3801 = _T_3799 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3290; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_3290[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3802 = _T_3801 & _GEN_634; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3795 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3797 = _T_3795 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3286; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_3286[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3798 = _T_3797 & _GEN_635; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3791 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3793 = _T_3791 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3282; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_3282[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3794 = _T_3793 & _GEN_636; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [599:0] _T_4289 = {_T_4280,_T_3826,_T_3822,_T_3818,_T_3814,_T_3810,_T_3806,_T_3802,_T_3798,_T_3794}; // @[Cat.scala 29:58]
  wire  _T_3787 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3789 = _T_3787 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3278; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_3278[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3790 = _T_3789 & _GEN_637; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3783 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3785 = _T_3783 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3274; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_3274[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3786 = _T_3785 & _GEN_638; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3779 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3781 = _T_3779 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3270; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_3270[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3782 = _T_3781 & _GEN_639; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3775 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3777 = _T_3775 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3266; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_3266[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3778 = _T_3777 & _GEN_640; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3771 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3773 = _T_3771 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3262; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_3262[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3774 = _T_3773 & _GEN_641; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3767 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3769 = _T_3767 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3258; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_3258[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3770 = _T_3769 & _GEN_642; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3763 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3765 = _T_3763 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3254; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_3254[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3766 = _T_3765 & _GEN_643; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3759 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3761 = _T_3759 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3250; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_3250[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3762 = _T_3761 & _GEN_644; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3755 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3757 = _T_3755 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3246; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_3246[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3758 = _T_3757 & _GEN_645; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [653:0] _T_4298 = {_T_4289,_T_3790,_T_3786,_T_3782,_T_3778,_T_3774,_T_3770,_T_3766,_T_3762,_T_3758}; // @[Cat.scala 29:58]
  wire  _T_3751 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3753 = _T_3751 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3242; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_3242[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3754 = _T_3753 & _GEN_646; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3747 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3749 = _T_3747 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3238; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_3238[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3750 = _T_3749 & _GEN_647; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3743 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3745 = _T_3743 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3234; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_3234[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3746 = _T_3745 & _GEN_648; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3739 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3741 = _T_3739 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3230; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_3230[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3742 = _T_3741 & _GEN_649; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3735 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3737 = _T_3735 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3226; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_3226[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3738 = _T_3737 & _GEN_650; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3731 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3733 = _T_3731 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3222; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_3222[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3734 = _T_3733 & _GEN_651; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3727 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3729 = _T_3727 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3218; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_3218[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3730 = _T_3729 & _GEN_652; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3723 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3725 = _T_3723 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3214; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_3214[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3726 = _T_3725 & _GEN_653; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3719 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3721 = _T_3719 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3210; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_3210[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3722 = _T_3721 & _GEN_654; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [707:0] _T_4307 = {_T_4298,_T_3754,_T_3750,_T_3746,_T_3742,_T_3738,_T_3734,_T_3730,_T_3726,_T_3722}; // @[Cat.scala 29:58]
  wire  _T_3715 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3717 = _T_3715 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3206; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_3206[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3718 = _T_3717 & _GEN_655; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3711 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3713 = _T_3711 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3202; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_3202[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3714 = _T_3713 & _GEN_656; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3707 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3709 = _T_3707 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3198; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_3198[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3710 = _T_3709 & _GEN_657; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3703 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3705 = _T_3703 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3194; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_3194[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3706 = _T_3705 & _GEN_658; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3699 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3701 = _T_3699 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3190; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_3190[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3702 = _T_3701 & _GEN_659; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3695 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3697 = _T_3695 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3186; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_3186[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3698 = _T_3697 & _GEN_660; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3691 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3693 = _T_3691 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3182; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_3182[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3694 = _T_3693 & _GEN_661; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3687 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3689 = _T_3687 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3178; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_3178[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3690 = _T_3689 & _GEN_662; // @[el2_ifu_mem_ctl.scala 729:130]
  wire  _T_3683 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3685 = _T_3683 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3174; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_3174[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3686 = _T_3685 & _GEN_663; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [761:0] _T_4316 = {_T_4307,_T_3718,_T_3714,_T_3710,_T_3706,_T_3702,_T_3698,_T_3694,_T_3690,_T_3686}; // @[Cat.scala 29:58]
  wire  _T_3679 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 729:121]
  wire [5:0] _T_3681 = _T_3679 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3170; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_3170[0]; // @[el2_ifu_mem_ctl.scala 726:30 el2_ifu_mem_ctl.scala 728:33]
  wire [5:0] _GEN_664 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [5:0] _T_3682 = _T_3681 & _GEN_664; // @[el2_ifu_mem_ctl.scala 729:130]
  wire [767:0] _T_4317 = {_T_4316,_T_3682}; // @[Cat.scala 29:58]
  wire  way_status = _T_4317[0]; // @[el2_ifu_mem_ctl.scala 729:16]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 262:96]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 264:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 266:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 271:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 276:59]
  wire  _T_214 = _T_212 | _T_1389; // @[el2_ifu_mem_ctl.scala 276:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 276:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 282:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 282:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 282:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 282:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 289:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 289:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 289:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 290:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 290:32]
  wire  _T_274 = imb_ff[12:6] == imb_scnd_ff[12:6]; // @[el2_ifu_mem_ctl.scala 293:75]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 293:127]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_1818 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 627:48]
  wire  _T_1819 = _T_1818 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 627:52]
  wire  bus_ifu_wr_data_error_ff = _T_1819 & miss_pending; // @[el2_ifu_mem_ctl.scala 627:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 372:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 371:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 293:145]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 293:143]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 296:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 296:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 297:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 316:30]
  wire  _T_9267 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 782:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 317:24]
  wire  _T_9269 = _T_9267 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 782:51]
  wire  _T_9271 = _T_9269 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 782:67]
  wire  _T_9273 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 782:86]
  wire  replace_way_mb_any_0 = _T_9271 | _T_9273; // @[el2_ifu_mem_ctl.scala 782:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9276 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 783:50]
  wire  _T_9278 = _T_9276 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 783:66]
  wire  _T_9280 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 783:85]
  wire  _T_9282 = _T_9280 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 783:100]
  wire  replace_way_mb_any_1 = _T_9278 | _T_9282; // @[el2_ifu_mem_ctl.scala 783:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 301:110]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 305:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 305:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 306:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 305:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 305:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 307:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 315:23]
  wire  _T_313 = _T_1404 & flush_final_f; // @[el2_ifu_mem_ctl.scala 319:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 319:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 319:53]
  wire  _T_1396 = ~_T_1391; // @[el2_ifu_mem_ctl.scala 462:46]
  wire  _T_1397 = _T_1389 & _T_1396; // @[el2_ifu_mem_ctl.scala 462:44]
  wire  stream_miss_f = _T_1397 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 462:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 319:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 319:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 325:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_1389; // @[el2_ifu_mem_ctl.scala 327:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 327:82]
  wire  _T_1410 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 467:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_1410}; // @[Cat.scala 29:58]
  wire  _T_1411 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 468:81]
  wire  _T_1435 = _T_1411 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1414 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 468:81]
  wire  _T_1436 = _T_1414 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1443 = _T_1435 | _T_1436; // @[Mux.scala 27:72]
  wire  _T_1417 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 468:81]
  wire  _T_1437 = _T_1417 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1444 = _T_1443 | _T_1437; // @[Mux.scala 27:72]
  wire  _T_1420 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 468:81]
  wire  _T_1438 = _T_1420 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1445 = _T_1444 | _T_1438; // @[Mux.scala 27:72]
  wire  _T_1423 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 468:81]
  wire  _T_1439 = _T_1423 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1445 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1426 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 468:81]
  wire  _T_1440 = _T_1426 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1429 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 468:81]
  wire  _T_1441 = _T_1429 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1432 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 468:81]
  wire  _T_1442 = _T_1432 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 469:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 331:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 331:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 624:61]
  wire  _T_1812 = ic_act_miss_f_delayed & _T_1405; // @[el2_ifu_mem_ctl.scala 625:53]
  wire  reset_tag_valid_for_miss = _T_1812 & _T_17; // @[el2_ifu_mem_ctl.scala 625:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 331:79]
  wire [30:0] _T_336 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_337 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 333:37]
  wire [30:0] _T_338 = sel_mb_addr ? _T_336 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_339 = _T_337 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_338 | _T_339; // @[Mux.scala 27:72]
  wire  _T_344 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 335:84]
  wire  _T_1806 = ~_T_1818; // @[el2_ifu_mem_ctl.scala 622:84]
  wire  _T_1807 = _T_100 & _T_1806; // @[el2_ifu_mem_ctl.scala 622:82]
  wire  bus_ifu_wr_en_ff_q = _T_1807 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 622:108]
  wire  sel_mb_status_addr = _T_344 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 335:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_336 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 336:31]
  wire [6:0] ic_wr_ecc = m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 345:13]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] ic_miss_buff_ecc = m2_io_ecc_out; // @[el2_ifu_mem_ctl.scala 348:20]
  wire [3:0] _T_1451 = {ifu_bus_rid_ff[2:1],_T_1410,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1452 = _T_1451 == 4'h0; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_1499 = _T_1452 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1455 = _T_1451 == 4'h1; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_1500 = _T_1455 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1515 = _T_1499 | _T_1500; // @[Mux.scala 27:72]
  wire  _T_1458 = _T_1451 == 4'h2; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_1501 = _T_1458 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1516 = _T_1515 | _T_1501; // @[Mux.scala 27:72]
  wire  _T_1461 = _T_1451 == 4'h3; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_1502 = _T_1461 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1517 = _T_1516 | _T_1502; // @[Mux.scala 27:72]
  wire  _T_1464 = _T_1451 == 4'h4; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_1503 = _T_1464 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1518 = _T_1517 | _T_1503; // @[Mux.scala 27:72]
  wire  _T_1467 = _T_1451 == 4'h5; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_1504 = _T_1467 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1519 = _T_1518 | _T_1504; // @[Mux.scala 27:72]
  wire  _T_1470 = _T_1451 == 4'h6; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_1505 = _T_1470 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1520 = _T_1519 | _T_1505; // @[Mux.scala 27:72]
  wire  _T_1473 = _T_1451 == 4'h7; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_1506 = _T_1473 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1521 = _T_1520 | _T_1506; // @[Mux.scala 27:72]
  wire  _T_1476 = _T_1451 == 4'h8; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_1507 = _T_1476 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1522 = _T_1521 | _T_1507; // @[Mux.scala 27:72]
  wire  _T_1479 = _T_1451 == 4'h9; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_1508 = _T_1479 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1523 = _T_1522 | _T_1508; // @[Mux.scala 27:72]
  wire  _T_1482 = _T_1451 == 4'ha; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_1509 = _T_1482 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1524 = _T_1523 | _T_1509; // @[Mux.scala 27:72]
  wire  _T_1485 = _T_1451 == 4'hb; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_1510 = _T_1485 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1525 = _T_1524 | _T_1510; // @[Mux.scala 27:72]
  wire  _T_1488 = _T_1451 == 4'hc; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_1511 = _T_1488 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1526 = _T_1525 | _T_1511; // @[Mux.scala 27:72]
  wire  _T_1491 = _T_1451 == 4'hd; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_1512 = _T_1491 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1527 = _T_1526 | _T_1512; // @[Mux.scala 27:72]
  wire  _T_1494 = _T_1451 == 4'he; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_1513 = _T_1494 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1528 = _T_1527 | _T_1513; // @[Mux.scala 27:72]
  wire  _T_1497 = _T_1451 == 4'hf; // @[el2_ifu_mem_ctl.scala 470:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_1514 = _T_1497 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1529 = _T_1528 | _T_1514; // @[Mux.scala 27:72]
  wire [3:0] _T_1531 = {ifu_bus_rid_ff[2:1],_T_1410,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1532 = _T_1531 == 4'h0; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1579 = _T_1532 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1535 = _T_1531 == 4'h1; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1580 = _T_1535 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1595 = _T_1579 | _T_1580; // @[Mux.scala 27:72]
  wire  _T_1538 = _T_1531 == 4'h2; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1581 = _T_1538 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1596 = _T_1595 | _T_1581; // @[Mux.scala 27:72]
  wire  _T_1541 = _T_1531 == 4'h3; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1582 = _T_1541 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1597 = _T_1596 | _T_1582; // @[Mux.scala 27:72]
  wire  _T_1544 = _T_1531 == 4'h4; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1583 = _T_1544 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1598 = _T_1597 | _T_1583; // @[Mux.scala 27:72]
  wire  _T_1547 = _T_1531 == 4'h5; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1584 = _T_1547 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1599 = _T_1598 | _T_1584; // @[Mux.scala 27:72]
  wire  _T_1550 = _T_1531 == 4'h6; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1585 = _T_1550 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1600 = _T_1599 | _T_1585; // @[Mux.scala 27:72]
  wire  _T_1553 = _T_1531 == 4'h7; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1586 = _T_1553 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1601 = _T_1600 | _T_1586; // @[Mux.scala 27:72]
  wire  _T_1556 = _T_1531 == 4'h8; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1587 = _T_1556 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1602 = _T_1601 | _T_1587; // @[Mux.scala 27:72]
  wire  _T_1559 = _T_1531 == 4'h9; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1588 = _T_1559 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1603 = _T_1602 | _T_1588; // @[Mux.scala 27:72]
  wire  _T_1562 = _T_1531 == 4'ha; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1589 = _T_1562 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1604 = _T_1603 | _T_1589; // @[Mux.scala 27:72]
  wire  _T_1565 = _T_1531 == 4'hb; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1590 = _T_1565 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1605 = _T_1604 | _T_1590; // @[Mux.scala 27:72]
  wire  _T_1568 = _T_1531 == 4'hc; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1591 = _T_1568 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1606 = _T_1605 | _T_1591; // @[Mux.scala 27:72]
  wire  _T_1571 = _T_1531 == 4'hd; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1592 = _T_1571 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1607 = _T_1606 | _T_1592; // @[Mux.scala 27:72]
  wire  _T_1574 = _T_1531 == 4'he; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1593 = _T_1574 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1608 = _T_1607 | _T_1593; // @[Mux.scala 27:72]
  wire  _T_1577 = _T_1531 == 4'hf; // @[el2_ifu_mem_ctl.scala 471:66]
  wire [31:0] _T_1594 = _T_1577 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1609 = _T_1608 | _T_1594; // @[Mux.scala 27:72]
  wire [141:0] _T_390 = {ic_wr_ecc,ifu_bus_rdata_ff,ic_miss_buff_ecc,_T_1529,_T_1609}; // @[Cat.scala 29:58]
  wire [141:0] _T_393 = {ic_miss_buff_ecc,_T_1529,_T_1609,ic_wr_ecc,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_390 : _T_393; // @[el2_ifu_mem_ctl.scala 363:28]
  wire  _T_352 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 353:56]
  wire  _T_353 = _T_352 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 353:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 417:28]
  wire  _T_569 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 419:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 620:35]
  wire  _T_438 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 402:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_438; // @[el2_ifu_mem_ctl.scala 402:73]
  wire  _T_495 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 408:118]
  wire  _T_496 = ic_miss_buff_data_valid[0] & _T_495; // @[el2_ifu_mem_ctl.scala 408:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_496; // @[el2_ifu_mem_ctl.scala 408:88]
  wire  _T_592 = _T_569 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_572 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 419:114]
  wire  _T_439 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 402:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_439; // @[el2_ifu_mem_ctl.scala 402:73]
  wire  _T_499 = ic_miss_buff_data_valid[1] & _T_495; // @[el2_ifu_mem_ctl.scala 408:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_499; // @[el2_ifu_mem_ctl.scala 408:88]
  wire  _T_593 = _T_572 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_600 = _T_592 | _T_593; // @[Mux.scala 27:72]
  wire  _T_575 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 419:114]
  wire  _T_440 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 402:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_440; // @[el2_ifu_mem_ctl.scala 402:73]
  wire  _T_502 = ic_miss_buff_data_valid[2] & _T_495; // @[el2_ifu_mem_ctl.scala 408:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_502; // @[el2_ifu_mem_ctl.scala 408:88]
  wire  _T_594 = _T_575 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_601 = _T_600 | _T_594; // @[Mux.scala 27:72]
  wire  _T_578 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 419:114]
  wire  _T_441 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 402:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_441; // @[el2_ifu_mem_ctl.scala 402:73]
  wire  _T_505 = ic_miss_buff_data_valid[3] & _T_495; // @[el2_ifu_mem_ctl.scala 408:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_505; // @[el2_ifu_mem_ctl.scala 408:88]
  wire  _T_595 = _T_578 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_602 = _T_601 | _T_595; // @[Mux.scala 27:72]
  wire  _T_581 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 419:114]
  wire  _T_442 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 402:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_442; // @[el2_ifu_mem_ctl.scala 402:73]
  wire  _T_508 = ic_miss_buff_data_valid[4] & _T_495; // @[el2_ifu_mem_ctl.scala 408:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_508; // @[el2_ifu_mem_ctl.scala 408:88]
  wire  _T_596 = _T_581 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_603 = _T_602 | _T_596; // @[Mux.scala 27:72]
  wire  _T_584 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 419:114]
  wire  _T_443 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 402:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_443; // @[el2_ifu_mem_ctl.scala 402:73]
  wire  _T_511 = ic_miss_buff_data_valid[5] & _T_495; // @[el2_ifu_mem_ctl.scala 408:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_511; // @[el2_ifu_mem_ctl.scala 408:88]
  wire  _T_597 = _T_584 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_604 = _T_603 | _T_597; // @[Mux.scala 27:72]
  wire  _T_587 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 419:114]
  wire  _T_444 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 402:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_444; // @[el2_ifu_mem_ctl.scala 402:73]
  wire  _T_514 = ic_miss_buff_data_valid[6] & _T_495; // @[el2_ifu_mem_ctl.scala 408:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_514; // @[el2_ifu_mem_ctl.scala 408:88]
  wire  _T_598 = _T_587 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_605 = _T_604 | _T_598; // @[Mux.scala 27:72]
  wire  _T_590 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 419:114]
  wire  _T_445 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 402:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_445; // @[el2_ifu_mem_ctl.scala 402:73]
  wire  _T_517 = ic_miss_buff_data_valid[7] & _T_495; // @[el2_ifu_mem_ctl.scala 408:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_517; // @[el2_ifu_mem_ctl.scala 408:88]
  wire  _T_599 = _T_590 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_605 | _T_599; // @[Mux.scala 27:72]
  wire  _T_608 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 420:58]
  wire  _T_609 = bypass_valid_value_check & _T_608; // @[el2_ifu_mem_ctl.scala 420:56]
  wire  _T_611 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 420:77]
  wire  _T_612 = _T_609 & _T_611; // @[el2_ifu_mem_ctl.scala 420:75]
  wire  _T_617 = _T_609 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 421:75]
  wire  _T_618 = _T_612 | _T_617; // @[el2_ifu_mem_ctl.scala 420:95]
  wire  _T_620 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 422:56]
  wire  _T_623 = _T_620 & _T_611; // @[el2_ifu_mem_ctl.scala 422:74]
  wire  _T_624 = _T_618 | _T_623; // @[el2_ifu_mem_ctl.scala 421:94]
  wire  _T_628 = _T_620 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 423:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 418:70]
  wire  _T_629 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 423:132]
  wire  _T_645 = _T_629 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_631 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 423:132]
  wire  _T_646 = _T_631 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_653 = _T_645 | _T_646; // @[Mux.scala 27:72]
  wire  _T_633 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 423:132]
  wire  _T_647 = _T_633 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_654 = _T_653 | _T_647; // @[Mux.scala 27:72]
  wire  _T_635 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 423:132]
  wire  _T_648 = _T_635 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_655 = _T_654 | _T_648; // @[Mux.scala 27:72]
  wire  _T_637 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 423:132]
  wire  _T_649 = _T_637 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_656 = _T_655 | _T_649; // @[Mux.scala 27:72]
  wire  _T_639 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 423:132]
  wire  _T_650 = _T_639 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_657 = _T_656 | _T_650; // @[Mux.scala 27:72]
  wire  _T_641 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 423:132]
  wire  _T_651 = _T_641 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_658 = _T_657 | _T_651; // @[Mux.scala 27:72]
  wire  _T_643 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 423:132]
  wire  _T_652 = _T_643 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_659 = _T_658 | _T_652; // @[Mux.scala 27:72]
  wire  _T_661 = _T_628 & _T_659; // @[el2_ifu_mem_ctl.scala 423:69]
  wire  _T_662 = _T_624 | _T_661; // @[el2_ifu_mem_ctl.scala 422:94]
  wire [4:0] _GEN_665 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 424:95]
  wire  _T_665 = _GEN_665 == 5'h1f; // @[el2_ifu_mem_ctl.scala 424:95]
  wire  _T_666 = bypass_valid_value_check & _T_665; // @[el2_ifu_mem_ctl.scala 424:56]
  wire  bypass_data_ready_in = _T_662 | _T_666; // @[el2_ifu_mem_ctl.scala 423:181]
  wire  _T_667 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 428:53]
  wire  _T_668 = _T_667 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 428:73]
  wire  _T_670 = _T_668 & _T_317; // @[el2_ifu_mem_ctl.scala 428:96]
  wire  _T_672 = _T_670 & _T_58; // @[el2_ifu_mem_ctl.scala 428:118]
  wire  _T_674 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 429:73]
  wire  _T_676 = _T_674 & _T_317; // @[el2_ifu_mem_ctl.scala 429:96]
  wire  _T_678 = _T_676 & _T_58; // @[el2_ifu_mem_ctl.scala 429:118]
  wire  _T_679 = _T_672 | _T_678; // @[el2_ifu_mem_ctl.scala 428:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 431:58]
  wire  _T_680 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 430:54]
  wire  _T_681 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 430:76]
  wire  _T_682 = _T_680 & _T_681; // @[el2_ifu_mem_ctl.scala 430:74]
  wire  _T_684 = _T_682 & _T_317; // @[el2_ifu_mem_ctl.scala 430:96]
  wire  ic_crit_wd_rdy_new_in = _T_679 | _T_684; // @[el2_ifu_mem_ctl.scala 429:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 630:43]
  wire  _T_405 = ic_crit_wd_rdy | _T_1389; // @[el2_ifu_mem_ctl.scala 376:38]
  wire  _T_407 = _T_405 | _T_1405; // @[el2_ifu_mem_ctl.scala 376:64]
  wire  _T_408 = ~_T_407; // @[el2_ifu_mem_ctl.scala 376:21]
  wire  _T_409 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 376:98]
  wire  sel_ic_data = _T_408 & _T_409; // @[el2_ifu_mem_ctl.scala 376:96]
  wire  _T_1612 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 475:44]
  wire  _T_778 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 442:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 414:60]
  wire  _T_722 = _T_569 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_723 = _T_572 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_730 = _T_722 | _T_723; // @[Mux.scala 27:72]
  wire  _T_724 = _T_575 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_731 = _T_730 | _T_724; // @[Mux.scala 27:72]
  wire  _T_725 = _T_578 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_732 = _T_731 | _T_725; // @[Mux.scala 27:72]
  wire  _T_726 = _T_581 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_733 = _T_732 | _T_726; // @[Mux.scala 27:72]
  wire  _T_727 = _T_584 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_734 = _T_733 | _T_727; // @[Mux.scala 27:72]
  wire  _T_728 = _T_587 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_735 = _T_734 | _T_728; // @[Mux.scala 27:72]
  wire  _T_729 = _T_590 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_735 | _T_729; // @[Mux.scala 27:72]
  wire  _T_761 = _T_1322 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_762 = _T_1325 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_769 = _T_761 | _T_762; // @[Mux.scala 27:72]
  wire  _T_763 = _T_1328 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_770 = _T_769 | _T_763; // @[Mux.scala 27:72]
  wire  _T_764 = _T_1331 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_771 = _T_770 | _T_764; // @[Mux.scala 27:72]
  wire  _T_765 = _T_1334 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_772 = _T_771 | _T_765; // @[Mux.scala 27:72]
  wire  _T_766 = _T_1337 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_773 = _T_772 | _T_766; // @[Mux.scala 27:72]
  wire  _T_767 = _T_1340 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_774 = _T_773 | _T_767; // @[Mux.scala 27:72]
  wire  _T_768 = _T_1343 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_774 | _T_768; // @[Mux.scala 27:72]
  wire  _T_779 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 444:70]
  wire  ifu_byp_data_err_new = _T_778 ? ic_miss_buff_data_error_bypass : _T_779; // @[el2_ifu_mem_ctl.scala 442:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 387:42]
  wire  _T_1613 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 475:91]
  wire  _T_1614 = ~_T_1613; // @[el2_ifu_mem_ctl.scala 475:60]
  wire  ic_rd_parity_final_err = _T_1612 & _T_1614; // @[el2_ifu_mem_ctl.scala 475:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_8885 = _T_3679 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 757:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_8887 = _T_3683 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9140 = _T_8885 | _T_8887; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_8889 = _T_3687 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9141 = _T_9140 | _T_8889; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_8891 = _T_3691 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9142 = _T_9141 | _T_8891; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_8893 = _T_3695 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9143 = _T_9142 | _T_8893; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_8895 = _T_3699 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9144 = _T_9143 | _T_8895; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_8897 = _T_3703 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9145 = _T_9144 | _T_8897; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_8899 = _T_3707 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9146 = _T_9145 | _T_8899; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_8901 = _T_3711 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9147 = _T_9146 | _T_8901; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_8903 = _T_3715 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9148 = _T_9147 | _T_8903; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_8905 = _T_3719 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9149 = _T_9148 | _T_8905; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_8907 = _T_3723 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9150 = _T_9149 | _T_8907; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_8909 = _T_3727 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9151 = _T_9150 | _T_8909; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_8911 = _T_3731 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9152 = _T_9151 | _T_8911; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_8913 = _T_3735 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9153 = _T_9152 | _T_8913; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_8915 = _T_3739 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9154 = _T_9153 | _T_8915; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_8917 = _T_3743 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9155 = _T_9154 | _T_8917; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_8919 = _T_3747 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9156 = _T_9155 | _T_8919; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_8921 = _T_3751 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9157 = _T_9156 | _T_8921; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_8923 = _T_3755 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9158 = _T_9157 | _T_8923; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_8925 = _T_3759 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9159 = _T_9158 | _T_8925; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_8927 = _T_3763 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9160 = _T_9159 | _T_8927; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_8929 = _T_3767 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9161 = _T_9160 | _T_8929; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_8931 = _T_3771 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9162 = _T_9161 | _T_8931; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_8933 = _T_3775 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9163 = _T_9162 | _T_8933; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_8935 = _T_3779 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9164 = _T_9163 | _T_8935; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_8937 = _T_3783 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9165 = _T_9164 | _T_8937; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_8939 = _T_3787 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9166 = _T_9165 | _T_8939; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_8941 = _T_3791 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9167 = _T_9166 | _T_8941; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_8943 = _T_3795 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9168 = _T_9167 | _T_8943; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_8945 = _T_3799 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9169 = _T_9168 | _T_8945; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_8947 = _T_3803 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9170 = _T_9169 | _T_8947; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_8949 = _T_3807 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9171 = _T_9170 | _T_8949; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_8951 = _T_3811 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9172 = _T_9171 | _T_8951; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_8953 = _T_3815 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9173 = _T_9172 | _T_8953; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_8955 = _T_3819 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9174 = _T_9173 | _T_8955; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_8957 = _T_3823 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9175 = _T_9174 | _T_8957; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_8959 = _T_3827 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9176 = _T_9175 | _T_8959; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_8961 = _T_3831 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9177 = _T_9176 | _T_8961; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_8963 = _T_3835 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9178 = _T_9177 | _T_8963; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_8965 = _T_3839 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9179 = _T_9178 | _T_8965; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_8967 = _T_3843 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9180 = _T_9179 | _T_8967; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_8969 = _T_3847 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9181 = _T_9180 | _T_8969; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_8971 = _T_3851 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9182 = _T_9181 | _T_8971; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_8973 = _T_3855 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9183 = _T_9182 | _T_8973; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_8975 = _T_3859 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9184 = _T_9183 | _T_8975; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_8977 = _T_3863 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9185 = _T_9184 | _T_8977; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_8979 = _T_3867 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9186 = _T_9185 | _T_8979; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_8981 = _T_3871 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9187 = _T_9186 | _T_8981; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_8983 = _T_3875 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9188 = _T_9187 | _T_8983; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_8985 = _T_3879 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9189 = _T_9188 | _T_8985; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_8987 = _T_3883 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9190 = _T_9189 | _T_8987; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_8989 = _T_3887 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9191 = _T_9190 | _T_8989; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_8991 = _T_3891 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9192 = _T_9191 | _T_8991; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_8993 = _T_3895 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9193 = _T_9192 | _T_8993; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_8995 = _T_3899 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9194 = _T_9193 | _T_8995; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_8997 = _T_3903 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9195 = _T_9194 | _T_8997; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_8999 = _T_3907 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9196 = _T_9195 | _T_8999; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9001 = _T_3911 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9197 = _T_9196 | _T_9001; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9003 = _T_3915 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9198 = _T_9197 | _T_9003; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9005 = _T_3919 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9199 = _T_9198 | _T_9005; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9007 = _T_3923 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9200 = _T_9199 | _T_9007; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9009 = _T_3927 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9201 = _T_9200 | _T_9009; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9011 = _T_3931 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9202 = _T_9201 | _T_9011; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9013 = _T_3935 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9203 = _T_9202 | _T_9013; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9015 = _T_3939 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9204 = _T_9203 | _T_9015; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9017 = _T_3943 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9205 = _T_9204 | _T_9017; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9019 = _T_3947 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9206 = _T_9205 | _T_9019; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9021 = _T_3951 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9207 = _T_9206 | _T_9021; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9023 = _T_3955 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9208 = _T_9207 | _T_9023; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9025 = _T_3959 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9209 = _T_9208 | _T_9025; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9027 = _T_3963 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9210 = _T_9209 | _T_9027; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9029 = _T_3967 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9211 = _T_9210 | _T_9029; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9031 = _T_3971 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9212 = _T_9211 | _T_9031; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9033 = _T_3975 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9213 = _T_9212 | _T_9033; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9035 = _T_3979 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9214 = _T_9213 | _T_9035; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9037 = _T_3983 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9215 = _T_9214 | _T_9037; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9039 = _T_3987 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9216 = _T_9215 | _T_9039; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9041 = _T_3991 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9217 = _T_9216 | _T_9041; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9043 = _T_3995 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9218 = _T_9217 | _T_9043; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9045 = _T_3999 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9219 = _T_9218 | _T_9045; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9047 = _T_4003 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9220 = _T_9219 | _T_9047; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9049 = _T_4007 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9221 = _T_9220 | _T_9049; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9051 = _T_4011 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9222 = _T_9221 | _T_9051; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9053 = _T_4015 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9223 = _T_9222 | _T_9053; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9055 = _T_4019 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9224 = _T_9223 | _T_9055; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9057 = _T_4023 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9225 = _T_9224 | _T_9057; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9059 = _T_4027 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9226 = _T_9225 | _T_9059; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9061 = _T_4031 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9227 = _T_9226 | _T_9061; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9063 = _T_4035 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9228 = _T_9227 | _T_9063; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9065 = _T_4039 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9229 = _T_9228 | _T_9065; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9067 = _T_4043 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9230 = _T_9229 | _T_9067; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9069 = _T_4047 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9231 = _T_9230 | _T_9069; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9071 = _T_4051 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9232 = _T_9231 | _T_9071; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9073 = _T_4055 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9233 = _T_9232 | _T_9073; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9075 = _T_4059 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9234 = _T_9233 | _T_9075; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9077 = _T_4063 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9235 = _T_9234 | _T_9077; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9079 = _T_4067 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9236 = _T_9235 | _T_9079; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9081 = _T_4071 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9237 = _T_9236 | _T_9081; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9083 = _T_4075 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9238 = _T_9237 | _T_9083; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9085 = _T_4079 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9239 = _T_9238 | _T_9085; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9087 = _T_4083 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9240 = _T_9239 | _T_9087; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9089 = _T_4087 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9241 = _T_9240 | _T_9089; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9091 = _T_4091 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9242 = _T_9241 | _T_9091; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9093 = _T_4095 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9243 = _T_9242 | _T_9093; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9095 = _T_4099 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9244 = _T_9243 | _T_9095; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9097 = _T_4103 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9245 = _T_9244 | _T_9097; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9099 = _T_4107 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9246 = _T_9245 | _T_9099; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9101 = _T_4111 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9247 = _T_9246 | _T_9101; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9103 = _T_4115 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9248 = _T_9247 | _T_9103; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9105 = _T_4119 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9249 = _T_9248 | _T_9105; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9107 = _T_4123 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9250 = _T_9249 | _T_9107; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9109 = _T_4127 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9251 = _T_9250 | _T_9109; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9111 = _T_4131 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9252 = _T_9251 | _T_9111; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9113 = _T_4135 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9253 = _T_9252 | _T_9113; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9115 = _T_4139 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9254 = _T_9253 | _T_9115; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9117 = _T_4143 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9255 = _T_9254 | _T_9117; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9119 = _T_4147 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9256 = _T_9255 | _T_9119; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9121 = _T_4151 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9257 = _T_9256 | _T_9121; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9123 = _T_4155 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9258 = _T_9257 | _T_9123; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9125 = _T_4159 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9259 = _T_9258 | _T_9125; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9127 = _T_4163 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9260 = _T_9259 | _T_9127; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9129 = _T_4167 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9261 = _T_9260 | _T_9129; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9131 = _T_4171 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9262 = _T_9261 | _T_9131; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9133 = _T_4175 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9263 = _T_9262 | _T_9133; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9135 = _T_4179 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9264 = _T_9263 | _T_9135; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9137 = _T_4183 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9265 = _T_9264 | _T_9137; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9139 = _T_4187 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_9266 = _T_9265 | _T_9139; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8502 = _T_3679 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 757:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8504 = _T_3683 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8757 = _T_8502 | _T_8504; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8506 = _T_3687 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8758 = _T_8757 | _T_8506; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8508 = _T_3691 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8759 = _T_8758 | _T_8508; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8510 = _T_3695 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8760 = _T_8759 | _T_8510; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_8512 = _T_3699 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8761 = _T_8760 | _T_8512; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_8514 = _T_3703 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8762 = _T_8761 | _T_8514; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_8516 = _T_3707 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8763 = _T_8762 | _T_8516; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_8518 = _T_3711 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8764 = _T_8763 | _T_8518; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_8520 = _T_3715 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8765 = _T_8764 | _T_8520; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_8522 = _T_3719 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8766 = _T_8765 | _T_8522; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_8524 = _T_3723 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8767 = _T_8766 | _T_8524; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_8526 = _T_3727 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8768 = _T_8767 | _T_8526; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_8528 = _T_3731 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8769 = _T_8768 | _T_8528; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_8530 = _T_3735 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8770 = _T_8769 | _T_8530; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_8532 = _T_3739 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8771 = _T_8770 | _T_8532; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_8534 = _T_3743 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8772 = _T_8771 | _T_8534; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_8536 = _T_3747 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8773 = _T_8772 | _T_8536; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_8538 = _T_3751 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8774 = _T_8773 | _T_8538; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_8540 = _T_3755 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8775 = _T_8774 | _T_8540; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_8542 = _T_3759 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8776 = _T_8775 | _T_8542; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_8544 = _T_3763 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8777 = _T_8776 | _T_8544; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_8546 = _T_3767 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8778 = _T_8777 | _T_8546; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_8548 = _T_3771 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8779 = _T_8778 | _T_8548; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_8550 = _T_3775 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8780 = _T_8779 | _T_8550; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_8552 = _T_3779 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8781 = _T_8780 | _T_8552; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_8554 = _T_3783 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8782 = _T_8781 | _T_8554; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_8556 = _T_3787 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8783 = _T_8782 | _T_8556; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_8558 = _T_3791 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8784 = _T_8783 | _T_8558; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_8560 = _T_3795 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8785 = _T_8784 | _T_8560; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_8562 = _T_3799 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8786 = _T_8785 | _T_8562; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_8564 = _T_3803 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8787 = _T_8786 | _T_8564; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_8566 = _T_3807 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8788 = _T_8787 | _T_8566; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_8568 = _T_3811 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8789 = _T_8788 | _T_8568; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_8570 = _T_3815 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8790 = _T_8789 | _T_8570; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_8572 = _T_3819 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8791 = _T_8790 | _T_8572; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_8574 = _T_3823 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8792 = _T_8791 | _T_8574; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_8576 = _T_3827 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8793 = _T_8792 | _T_8576; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_8578 = _T_3831 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8794 = _T_8793 | _T_8578; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_8580 = _T_3835 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8795 = _T_8794 | _T_8580; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_8582 = _T_3839 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8796 = _T_8795 | _T_8582; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_8584 = _T_3843 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8797 = _T_8796 | _T_8584; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_8586 = _T_3847 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8798 = _T_8797 | _T_8586; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_8588 = _T_3851 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8799 = _T_8798 | _T_8588; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_8590 = _T_3855 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8800 = _T_8799 | _T_8590; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_8592 = _T_3859 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8801 = _T_8800 | _T_8592; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_8594 = _T_3863 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8802 = _T_8801 | _T_8594; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_8596 = _T_3867 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8803 = _T_8802 | _T_8596; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_8598 = _T_3871 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8804 = _T_8803 | _T_8598; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_8600 = _T_3875 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8805 = _T_8804 | _T_8600; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_8602 = _T_3879 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8806 = _T_8805 | _T_8602; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_8604 = _T_3883 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8807 = _T_8806 | _T_8604; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_8606 = _T_3887 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8808 = _T_8807 | _T_8606; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_8608 = _T_3891 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8809 = _T_8808 | _T_8608; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_8610 = _T_3895 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8810 = _T_8809 | _T_8610; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_8612 = _T_3899 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8811 = _T_8810 | _T_8612; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_8614 = _T_3903 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8812 = _T_8811 | _T_8614; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_8616 = _T_3907 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8813 = _T_8812 | _T_8616; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_8618 = _T_3911 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8814 = _T_8813 | _T_8618; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_8620 = _T_3915 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8815 = _T_8814 | _T_8620; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_8622 = _T_3919 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8816 = _T_8815 | _T_8622; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_8624 = _T_3923 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8817 = _T_8816 | _T_8624; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_8626 = _T_3927 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8818 = _T_8817 | _T_8626; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_8628 = _T_3931 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8819 = _T_8818 | _T_8628; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_8630 = _T_3935 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8820 = _T_8819 | _T_8630; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_8632 = _T_3939 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8821 = _T_8820 | _T_8632; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_8634 = _T_3943 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8822 = _T_8821 | _T_8634; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_8636 = _T_3947 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8823 = _T_8822 | _T_8636; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_8638 = _T_3951 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8824 = _T_8823 | _T_8638; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_8640 = _T_3955 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8825 = _T_8824 | _T_8640; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_8642 = _T_3959 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8826 = _T_8825 | _T_8642; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_8644 = _T_3963 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8827 = _T_8826 | _T_8644; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_8646 = _T_3967 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8828 = _T_8827 | _T_8646; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_8648 = _T_3971 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8829 = _T_8828 | _T_8648; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_8650 = _T_3975 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8830 = _T_8829 | _T_8650; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_8652 = _T_3979 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8831 = _T_8830 | _T_8652; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_8654 = _T_3983 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8832 = _T_8831 | _T_8654; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_8656 = _T_3987 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8833 = _T_8832 | _T_8656; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_8658 = _T_3991 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8834 = _T_8833 | _T_8658; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_8660 = _T_3995 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8835 = _T_8834 | _T_8660; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_8662 = _T_3999 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8836 = _T_8835 | _T_8662; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_8664 = _T_4003 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8837 = _T_8836 | _T_8664; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_8666 = _T_4007 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8838 = _T_8837 | _T_8666; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_8668 = _T_4011 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8839 = _T_8838 | _T_8668; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_8670 = _T_4015 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8840 = _T_8839 | _T_8670; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_8672 = _T_4019 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8841 = _T_8840 | _T_8672; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_8674 = _T_4023 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8842 = _T_8841 | _T_8674; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_8676 = _T_4027 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8843 = _T_8842 | _T_8676; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_8678 = _T_4031 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8844 = _T_8843 | _T_8678; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_8680 = _T_4035 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8845 = _T_8844 | _T_8680; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_8682 = _T_4039 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8846 = _T_8845 | _T_8682; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_8684 = _T_4043 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8847 = _T_8846 | _T_8684; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_8686 = _T_4047 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8848 = _T_8847 | _T_8686; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_8688 = _T_4051 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8849 = _T_8848 | _T_8688; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_8690 = _T_4055 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8850 = _T_8849 | _T_8690; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_8692 = _T_4059 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8851 = _T_8850 | _T_8692; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_8694 = _T_4063 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8852 = _T_8851 | _T_8694; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_8696 = _T_4067 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8853 = _T_8852 | _T_8696; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_8698 = _T_4071 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8854 = _T_8853 | _T_8698; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_8700 = _T_4075 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8855 = _T_8854 | _T_8700; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_8702 = _T_4079 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8856 = _T_8855 | _T_8702; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_8704 = _T_4083 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8857 = _T_8856 | _T_8704; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_8706 = _T_4087 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8858 = _T_8857 | _T_8706; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_8708 = _T_4091 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8859 = _T_8858 | _T_8708; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_8710 = _T_4095 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8860 = _T_8859 | _T_8710; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_8712 = _T_4099 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8861 = _T_8860 | _T_8712; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_8714 = _T_4103 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8862 = _T_8861 | _T_8714; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_8716 = _T_4107 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8863 = _T_8862 | _T_8716; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_8718 = _T_4111 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8864 = _T_8863 | _T_8718; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_8720 = _T_4115 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8865 = _T_8864 | _T_8720; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_8722 = _T_4119 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8866 = _T_8865 | _T_8722; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_8724 = _T_4123 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8867 = _T_8866 | _T_8724; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_8726 = _T_4127 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8868 = _T_8867 | _T_8726; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_8728 = _T_4131 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8869 = _T_8868 | _T_8728; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_8730 = _T_4135 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8870 = _T_8869 | _T_8730; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_8732 = _T_4139 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8871 = _T_8870 | _T_8732; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_8734 = _T_4143 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8872 = _T_8871 | _T_8734; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_8736 = _T_4147 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8873 = _T_8872 | _T_8736; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_8738 = _T_4151 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8874 = _T_8873 | _T_8738; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_8740 = _T_4155 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8875 = _T_8874 | _T_8740; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_8742 = _T_4159 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8876 = _T_8875 | _T_8742; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_8744 = _T_4163 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8877 = _T_8876 | _T_8744; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_8746 = _T_4167 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8878 = _T_8877 | _T_8746; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_8748 = _T_4171 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8879 = _T_8878 | _T_8748; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_8750 = _T_4175 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8880 = _T_8879 | _T_8750; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_8752 = _T_4179 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8881 = _T_8880 | _T_8752; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_8754 = _T_4183 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8882 = _T_8881 | _T_8754; // @[el2_ifu_mem_ctl.scala 757:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_8756 = _T_4187 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 757:10]
  wire  _T_8883 = _T_8882 | _T_8756; // @[el2_ifu_mem_ctl.scala 757:91]
  wire [1:0] ic_tag_valid_unq = {_T_9266,_T_8883}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 830:54]
  wire [1:0] _T_9305 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9306 = ic_debug_way_ff & _T_9305; // @[el2_ifu_mem_ctl.scala 811:67]
  wire [1:0] _T_9307 = ic_tag_valid_unq & _T_9306; // @[el2_ifu_mem_ctl.scala 811:48]
  wire  ic_debug_tag_val_rd_out = |_T_9307; // @[el2_ifu_mem_ctl.scala 811:115]
  wire [65:0] _T_364 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_365; // @[Reg.scala 27:20]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_1747; // @[el2_ifu_mem_ctl.scala 370:80]
  wire  _T_403 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 375:98]
  wire  sel_byp_data = _T_407 & _T_403; // @[el2_ifu_mem_ctl.scala 375:96]
  wire [63:0] _T_414 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_415 = _T_414 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 382:64]
  wire [63:0] _T_417 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_1269 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 450:31]
  wire  _T_782 = ~ifu_fetch_addr_int_f[1]; // @[el2_ifu_mem_ctl.scala 446:38]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_783 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_831 = _T_783 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_786 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_832 = _T_786 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_847 = _T_831 | _T_832; // @[Mux.scala 27:72]
  wire  _T_789 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_833 = _T_789 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_848 = _T_847 | _T_833; // @[Mux.scala 27:72]
  wire  _T_792 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_834 = _T_792 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_849 = _T_848 | _T_834; // @[Mux.scala 27:72]
  wire  _T_795 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_835 = _T_795 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_850 = _T_849 | _T_835; // @[Mux.scala 27:72]
  wire  _T_798 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_836 = _T_798 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_851 = _T_850 | _T_836; // @[Mux.scala 27:72]
  wire  _T_801 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_837 = _T_801 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_852 = _T_851 | _T_837; // @[Mux.scala 27:72]
  wire  _T_804 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_838 = _T_804 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_853 = _T_852 | _T_838; // @[Mux.scala 27:72]
  wire  _T_807 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_839 = _T_807 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_854 = _T_853 | _T_839; // @[Mux.scala 27:72]
  wire  _T_810 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_840 = _T_810 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_855 = _T_854 | _T_840; // @[Mux.scala 27:72]
  wire  _T_813 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_841 = _T_813 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_856 = _T_855 | _T_841; // @[Mux.scala 27:72]
  wire  _T_816 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_842 = _T_816 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_857 = _T_856 | _T_842; // @[Mux.scala 27:72]
  wire  _T_819 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_843 = _T_819 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_858 = _T_857 | _T_843; // @[Mux.scala 27:72]
  wire  _T_822 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_844 = _T_822 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_859 = _T_858 | _T_844; // @[Mux.scala 27:72]
  wire  _T_825 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_845 = _T_825 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_860 = _T_859 | _T_845; // @[Mux.scala 27:72]
  wire  _T_828 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_846 = _T_828 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_861 = _T_860 | _T_846; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_863 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_911 = _T_863 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_866 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_912 = _T_866 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_927 = _T_911 | _T_912; // @[Mux.scala 27:72]
  wire  _T_869 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_913 = _T_869 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_928 = _T_927 | _T_913; // @[Mux.scala 27:72]
  wire  _T_872 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_914 = _T_872 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_929 = _T_928 | _T_914; // @[Mux.scala 27:72]
  wire  _T_875 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_915 = _T_875 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_930 = _T_929 | _T_915; // @[Mux.scala 27:72]
  wire  _T_878 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_916 = _T_878 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_931 = _T_930 | _T_916; // @[Mux.scala 27:72]
  wire  _T_881 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_917 = _T_881 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_932 = _T_931 | _T_917; // @[Mux.scala 27:72]
  wire  _T_884 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_918 = _T_884 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_933 = _T_932 | _T_918; // @[Mux.scala 27:72]
  wire  _T_887 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_919 = _T_887 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_934 = _T_933 | _T_919; // @[Mux.scala 27:72]
  wire  _T_890 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_920 = _T_890 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_935 = _T_934 | _T_920; // @[Mux.scala 27:72]
  wire  _T_893 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_921 = _T_893 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_936 = _T_935 | _T_921; // @[Mux.scala 27:72]
  wire  _T_896 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_922 = _T_896 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_937 = _T_936 | _T_922; // @[Mux.scala 27:72]
  wire  _T_899 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_923 = _T_899 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_938 = _T_937 | _T_923; // @[Mux.scala 27:72]
  wire  _T_902 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_924 = _T_902 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_939 = _T_938 | _T_924; // @[Mux.scala 27:72]
  wire  _T_905 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_925 = _T_905 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_940 = _T_939 | _T_925; // @[Mux.scala 27:72]
  wire  _T_908 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 447:179]
  wire [31:0] _T_926 = _T_908 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_941 = _T_940 | _T_926; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_943 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_991 = _T_943 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_946 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_992 = _T_946 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1007 = _T_991 | _T_992; // @[Mux.scala 27:72]
  wire  _T_949 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_993 = _T_949 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1008 = _T_1007 | _T_993; // @[Mux.scala 27:72]
  wire  _T_952 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_994 = _T_952 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1009 = _T_1008 | _T_994; // @[Mux.scala 27:72]
  wire  _T_955 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_995 = _T_955 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1010 = _T_1009 | _T_995; // @[Mux.scala 27:72]
  wire  _T_958 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_996 = _T_958 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1011 = _T_1010 | _T_996; // @[Mux.scala 27:72]
  wire  _T_961 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_997 = _T_961 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1012 = _T_1011 | _T_997; // @[Mux.scala 27:72]
  wire  _T_964 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_998 = _T_964 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1013 = _T_1012 | _T_998; // @[Mux.scala 27:72]
  wire  _T_967 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_999 = _T_967 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1014 = _T_1013 | _T_999; // @[Mux.scala 27:72]
  wire  _T_970 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_1000 = _T_970 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1015 = _T_1014 | _T_1000; // @[Mux.scala 27:72]
  wire  _T_973 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_1001 = _T_973 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1016 = _T_1015 | _T_1001; // @[Mux.scala 27:72]
  wire  _T_976 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_1002 = _T_976 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1017 = _T_1016 | _T_1002; // @[Mux.scala 27:72]
  wire  _T_979 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_1003 = _T_979 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1018 = _T_1017 | _T_1003; // @[Mux.scala 27:72]
  wire  _T_982 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_1004 = _T_982 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1019 = _T_1018 | _T_1004; // @[Mux.scala 27:72]
  wire  _T_985 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_1005 = _T_985 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1020 = _T_1019 | _T_1005; // @[Mux.scala 27:72]
  wire  _T_988 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 447:285]
  wire [31:0] _T_1006 = _T_988 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1021 = _T_1020 | _T_1006; // @[Mux.scala 27:72]
  wire [79:0] _T_1024 = {_T_861,_T_941,_T_1021}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1025 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1073 = _T_1025 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1028 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1074 = _T_1028 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1089 = _T_1073 | _T_1074; // @[Mux.scala 27:72]
  wire  _T_1031 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1075 = _T_1031 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1090 = _T_1089 | _T_1075; // @[Mux.scala 27:72]
  wire  _T_1034 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1076 = _T_1034 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1091 = _T_1090 | _T_1076; // @[Mux.scala 27:72]
  wire  _T_1037 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1077 = _T_1037 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1092 = _T_1091 | _T_1077; // @[Mux.scala 27:72]
  wire  _T_1040 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1078 = _T_1040 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1093 = _T_1092 | _T_1078; // @[Mux.scala 27:72]
  wire  _T_1043 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1079 = _T_1043 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1094 = _T_1093 | _T_1079; // @[Mux.scala 27:72]
  wire  _T_1046 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1080 = _T_1046 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1095 = _T_1094 | _T_1080; // @[Mux.scala 27:72]
  wire  _T_1049 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1081 = _T_1049 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1096 = _T_1095 | _T_1081; // @[Mux.scala 27:72]
  wire  _T_1052 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1082 = _T_1052 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1097 = _T_1096 | _T_1082; // @[Mux.scala 27:72]
  wire  _T_1055 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1083 = _T_1055 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1098 = _T_1097 | _T_1083; // @[Mux.scala 27:72]
  wire  _T_1058 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1084 = _T_1058 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1099 = _T_1098 | _T_1084; // @[Mux.scala 27:72]
  wire  _T_1061 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1085 = _T_1061 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1100 = _T_1099 | _T_1085; // @[Mux.scala 27:72]
  wire  _T_1064 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1086 = _T_1064 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1101 = _T_1100 | _T_1086; // @[Mux.scala 27:72]
  wire  _T_1067 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1087 = _T_1067 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1102 = _T_1101 | _T_1087; // @[Mux.scala 27:72]
  wire  _T_1070 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 448:73]
  wire [15:0] _T_1088 = _T_1070 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1103 = _T_1102 | _T_1088; // @[Mux.scala 27:72]
  wire [31:0] _T_1153 = _T_783 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1154 = _T_786 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1169 = _T_1153 | _T_1154; // @[Mux.scala 27:72]
  wire [31:0] _T_1155 = _T_789 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1170 = _T_1169 | _T_1155; // @[Mux.scala 27:72]
  wire [31:0] _T_1156 = _T_792 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1171 = _T_1170 | _T_1156; // @[Mux.scala 27:72]
  wire [31:0] _T_1157 = _T_795 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1172 = _T_1171 | _T_1157; // @[Mux.scala 27:72]
  wire [31:0] _T_1158 = _T_798 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1173 = _T_1172 | _T_1158; // @[Mux.scala 27:72]
  wire [31:0] _T_1159 = _T_801 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1174 = _T_1173 | _T_1159; // @[Mux.scala 27:72]
  wire [31:0] _T_1160 = _T_804 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1175 = _T_1174 | _T_1160; // @[Mux.scala 27:72]
  wire [31:0] _T_1161 = _T_807 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1176 = _T_1175 | _T_1161; // @[Mux.scala 27:72]
  wire [31:0] _T_1162 = _T_810 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1177 = _T_1176 | _T_1162; // @[Mux.scala 27:72]
  wire [31:0] _T_1163 = _T_813 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1178 = _T_1177 | _T_1163; // @[Mux.scala 27:72]
  wire [31:0] _T_1164 = _T_816 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1179 = _T_1178 | _T_1164; // @[Mux.scala 27:72]
  wire [31:0] _T_1165 = _T_819 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1180 = _T_1179 | _T_1165; // @[Mux.scala 27:72]
  wire [31:0] _T_1166 = _T_822 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1181 = _T_1180 | _T_1166; // @[Mux.scala 27:72]
  wire [31:0] _T_1167 = _T_825 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1182 = _T_1181 | _T_1167; // @[Mux.scala 27:72]
  wire [31:0] _T_1168 = _T_828 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1183 = _T_1182 | _T_1168; // @[Mux.scala 27:72]
  wire [79:0] _T_1266 = {_T_1103,_T_1183,_T_941}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_782 ? _T_1024 : _T_1266; // @[el2_ifu_mem_ctl.scala 446:37]
  wire [79:0] _T_1271 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_1269 ? ic_byp_data_only_pre_new : _T_1271; // @[el2_ifu_mem_ctl.scala 450:30]
  wire [79:0] _GEN_794 = {{16'd0}, _T_417}; // @[el2_ifu_mem_ctl.scala 382:109]
  wire [79:0] _T_418 = _GEN_794 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 382:109]
  wire [79:0] _GEN_795 = {{16'd0}, _T_415}; // @[el2_ifu_mem_ctl.scala 382:83]
  wire [79:0] ic_premux_data = _GEN_795 | _T_418; // @[el2_ifu_mem_ctl.scala 382:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 389:38]
  wire [1:0] _T_427 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 393:8]
  wire  _T_429 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[el2_ifu_mem_ctl.scala 395:45]
  wire  _T_431 = byp_fetch_index == 5'h1f; // @[el2_ifu_mem_ctl.scala 395:80]
  wire  _T_432 = ~_T_431; // @[el2_ifu_mem_ctl.scala 395:71]
  wire  _T_433 = _T_429 & _T_432; // @[el2_ifu_mem_ctl.scala 395:69]
  wire  _T_434 = err_stop_state != 2'h2; // @[el2_ifu_mem_ctl.scala 395:131]
  wire  _T_435 = _T_433 & _T_434; // @[el2_ifu_mem_ctl.scala 395:114]
  wire [7:0] _T_524 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_529 = ic_miss_buff_data_error[0] & _T_495; // @[el2_ifu_mem_ctl.scala 413:32]
  wire  _T_1815 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 626:47]
  wire  _T_1816 = _T_1815 & _T_13; // @[el2_ifu_mem_ctl.scala 626:50]
  wire  bus_ifu_wr_data_error = _T_1816 & miss_pending; // @[el2_ifu_mem_ctl.scala 626:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_529; // @[el2_ifu_mem_ctl.scala 412:72]
  wire  _T_533 = ic_miss_buff_data_error[1] & _T_495; // @[el2_ifu_mem_ctl.scala 413:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_533; // @[el2_ifu_mem_ctl.scala 412:72]
  wire  _T_537 = ic_miss_buff_data_error[2] & _T_495; // @[el2_ifu_mem_ctl.scala 413:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_537; // @[el2_ifu_mem_ctl.scala 412:72]
  wire  _T_541 = ic_miss_buff_data_error[3] & _T_495; // @[el2_ifu_mem_ctl.scala 413:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_541; // @[el2_ifu_mem_ctl.scala 412:72]
  wire  _T_545 = ic_miss_buff_data_error[4] & _T_495; // @[el2_ifu_mem_ctl.scala 413:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_545; // @[el2_ifu_mem_ctl.scala 412:72]
  wire  _T_549 = ic_miss_buff_data_error[5] & _T_495; // @[el2_ifu_mem_ctl.scala 413:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_549; // @[el2_ifu_mem_ctl.scala 412:72]
  wire  _T_553 = ic_miss_buff_data_error[6] & _T_495; // @[el2_ifu_mem_ctl.scala 413:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_553; // @[el2_ifu_mem_ctl.scala 412:72]
  wire  _T_557 = ic_miss_buff_data_error[7] & _T_495; // @[el2_ifu_mem_ctl.scala 413:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_557; // @[el2_ifu_mem_ctl.scala 412:72]
  wire [7:0] _T_564 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_1621 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1629 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 495:65]
  wire  _T_1630 = _T_1629 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 495:88]
  wire  _T_1632 = _T_1630 & _T_1743; // @[el2_ifu_mem_ctl.scala 495:112]
  wire  _T_1633 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1634 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 500:50]
  wire  _T_1636 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1642 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1644 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_39 = _T_1642 | _T_1644; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_1636 ? _T_1634 : _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_1633 ? _T_1634 : _GEN_41; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_1621 ? _T_1632 : _GEN_43; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_1621 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_1635 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 501:56]
  wire  _GEN_44 = _T_1633 & _T_1635; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_1621 ? 1'h0 : _GEN_44; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 486:58]
  wire  _T_1618 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 485:49]
  wire  _T_1623 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 494:87]
  wire  _T_1637 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 504:54]
  wire  _T_1638 = _T_1637 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 504:84]
  wire  _T_1647 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 525:66]
  wire  _T_1648 = io_dec_tlu_flush_err_wb & _T_1647; // @[el2_ifu_mem_ctl.scala 525:52]
  wire  _T_1650 = _T_1648 & _T_1743; // @[el2_ifu_mem_ctl.scala 525:81]
  wire  _T_1652 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 528:59]
  wire  _T_1653 = _T_1652 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 528:86]
  wire  _T_1667 = _T_1652 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 531:81]
  wire  _T_1668 = _T_1667 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 531:103]
  wire  _T_1669 = _T_1668 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 531:126]
  wire  _T_1689 = _T_1667 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 538:103]
  wire  _T_1696 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 543:62]
  wire  _T_1697 = io_dec_tlu_flush_lower_wb & _T_1696; // @[el2_ifu_mem_ctl.scala 543:60]
  wire  _T_1698 = _T_1697 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 543:88]
  wire  _T_1699 = _T_1698 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 543:115]
  wire  _GEN_51 = _T_1695 & _T_1653; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_1678 ? _T_1689 : _GEN_51; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_1678 | _T_1695; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_1651 ? _T_1669 : _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_1651 | _GEN_56; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_1646 ? _T_1650 : _GEN_58; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_1711 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 560:64]
  wire  _T_1713 = _T_1711 & _T_1743; // @[el2_ifu_mem_ctl.scala 560:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_1715 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 560:133]
  wire  _T_1716 = _T_1715 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 560:164]
  wire  _T_1717 = _T_1716 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 560:184]
  wire  _T_1718 = _T_1717 & miss_pending; // @[el2_ifu_mem_ctl.scala 560:204]
  wire  _T_1719 = ~_T_1718; // @[el2_ifu_mem_ctl.scala 560:112]
  wire  ifc_bus_ic_req_ff_in = _T_1713 & _T_1719; // @[el2_ifu_mem_ctl.scala 560:110]
  wire  _T_1720 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 561:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 592:45]
  wire  _T_1737 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 595:35]
  wire  _T_1738 = _T_1737 & miss_pending; // @[el2_ifu_mem_ctl.scala 595:53]
  wire  bus_cmd_sent = _T_1738 & _T_1743; // @[el2_ifu_mem_ctl.scala 595:68]
  wire [2:0] _T_1728 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1730 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_1732 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 593:51]
  wire  _T_1758 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 603:73]
  wire  _T_1759 = _T_1744 & _T_1758; // @[el2_ifu_mem_ctl.scala 603:71]
  wire  _T_1761 = last_data_recieved_ff & _T_495; // @[el2_ifu_mem_ctl.scala 603:114]
  wire  last_data_recieved_in = _T_1759 | _T_1761; // @[el2_ifu_mem_ctl.scala 603:89]
  wire [2:0] _T_1767 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 608:45]
  wire  _T_1770 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 609:81]
  wire  _T_1771 = _T_1770 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 609:97]
  wire  _T_1773 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 611:48]
  wire  _T_1774 = _T_1773 & miss_pending; // @[el2_ifu_mem_ctl.scala 611:68]
  wire  bus_inc_cmd_beat_cnt = _T_1774 & _T_1743; // @[el2_ifu_mem_ctl.scala 611:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 613:57]
  wire  _T_1778 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 614:31]
  wire  _T_1779 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 614:71]
  wire  _T_1780 = _T_1779 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 614:87]
  wire  _T_1781 = ~_T_1780; // @[el2_ifu_mem_ctl.scala 614:55]
  wire  bus_hold_cmd_beat_cnt = _T_1778 & _T_1781; // @[el2_ifu_mem_ctl.scala 614:53]
  wire  _T_1782 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 615:46]
  wire  bus_cmd_beat_en = _T_1782 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 615:62]
  wire [2:0] _T_1785 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 617:46]
  wire [2:0] _T_1787 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1788 = bus_inc_cmd_beat_cnt ? _T_1785 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1789 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1791 = _T_1787 | _T_1788; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_1791 | _T_1789; // @[Mux.scala 27:72]
  wire  _T_1795 = _T_1771 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 618:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 629:62]
  wire  _T_1823 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 634:50]
  wire  _T_1824 = io_ifc_dma_access_ok & _T_1823; // @[el2_ifu_mem_ctl.scala 634:47]
  wire  _T_1825 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 634:70]
  wire  ifc_dma_access_ok_d = _T_1824 & _T_1825; // @[el2_ifu_mem_ctl.scala 634:68]
  wire  _T_1829 = _T_1824 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 635:72]
  wire  _T_1830 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 635:111]
  wire  _T_1831 = _T_1829 & _T_1830; // @[el2_ifu_mem_ctl.scala 635:97]
  wire  ifc_dma_access_q_ok = _T_1831 & _T_1825; // @[el2_ifu_mem_ctl.scala 635:127]
  wire  _T_1834 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 638:40]
  wire  _T_1835 = _T_1834 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 638:58]
  wire  _T_1838 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 639:60]
  wire  _T_1839 = _T_1834 & _T_1838; // @[el2_ifu_mem_ctl.scala 639:58]
  wire  _T_1840 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 639:104]
  wire [2:0] _T_1845 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_1951 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_1960 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_1951}; // @[el2_lib.scala 268:22]
  wire  _T_1961 = ^_T_1960; // @[el2_lib.scala 268:29]
  wire [8:0] _T_1969 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_1978 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_1969}; // @[el2_lib.scala 268:39]
  wire  _T_1979 = ^_T_1978; // @[el2_lib.scala 268:46]
  wire [8:0] _T_1987 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_1996 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_1987}; // @[el2_lib.scala 268:56]
  wire  _T_1997 = ^_T_1996; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2003 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2011 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_2003}; // @[el2_lib.scala 268:73]
  wire  _T_2012 = ^_T_2011; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2026 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_2003}; // @[el2_lib.scala 268:90]
  wire  _T_2027 = ^_T_2026; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2032 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_2033 = ^_T_2032; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2038 = {_T_1961,_T_1979,_T_1997,_T_2012,_T_2027,_T_2033}; // @[Cat.scala 29:58]
  wire  _T_2039 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2040 = ^_T_2038; // @[el2_lib.scala 269:23]
  wire  _T_2041 = _T_2039 ^ _T_2040; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2147 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2156 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2147}; // @[el2_lib.scala 268:22]
  wire  _T_2157 = ^_T_2156; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2165 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2174 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_2165}; // @[el2_lib.scala 268:39]
  wire  _T_2175 = ^_T_2174; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2183 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2192 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_2183}; // @[el2_lib.scala 268:56]
  wire  _T_2193 = ^_T_2192; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2199 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2207 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_2199}; // @[el2_lib.scala 268:73]
  wire  _T_2208 = ^_T_2207; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2222 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_2199}; // @[el2_lib.scala 268:90]
  wire  _T_2223 = ^_T_2222; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2228 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_2229 = ^_T_2228; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2234 = {_T_2157,_T_2175,_T_2193,_T_2208,_T_2223,_T_2229}; // @[Cat.scala 29:58]
  wire  _T_2235 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_2236 = ^_T_2234; // @[el2_lib.scala 269:23]
  wire  _T_2237 = _T_2235 ^ _T_2236; // @[el2_lib.scala 269:18]
  wire [6:0] _T_2238 = {_T_2237,_T_2157,_T_2175,_T_2193,_T_2208,_T_2223,_T_2229}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2041,_T_1961,_T_1979,_T_1997,_T_2012,_T_2027,_T_2033,_T_2238}; // @[Cat.scala 29:58]
  wire  _T_2240 = ~_T_1834; // @[el2_ifu_mem_ctl.scala 644:45]
  wire  _T_2241 = iccm_correct_ecc & _T_2240; // @[el2_ifu_mem_ctl.scala 644:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_2242 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_2249 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 658:53]
  wire  _T_2581 = _T_2493[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_2579 = _T_2493[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_2577 = _T_2493[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_2575 = _T_2493[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_2573 = _T_2493[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_2571 = _T_2493[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_2569 = _T_2493[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_2567 = _T_2493[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_2565 = _T_2493[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_2563 = _T_2493[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2639 = {_T_2581,_T_2579,_T_2577,_T_2575,_T_2573,_T_2571,_T_2569,_T_2567,_T_2565,_T_2563}; // @[el2_lib.scala 310:69]
  wire  _T_2561 = _T_2493[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_2559 = _T_2493[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_2557 = _T_2493[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_2555 = _T_2493[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_2553 = _T_2493[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_2551 = _T_2493[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_2549 = _T_2493[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_2547 = _T_2493[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_2545 = _T_2493[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_2543 = _T_2493[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2630 = {_T_2561,_T_2559,_T_2557,_T_2555,_T_2553,_T_2551,_T_2549,_T_2547,_T_2545,_T_2543}; // @[el2_lib.scala 310:69]
  wire  _T_2541 = _T_2493[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_2539 = _T_2493[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_2537 = _T_2493[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_2535 = _T_2493[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_2533 = _T_2493[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_2531 = _T_2493[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_2529 = _T_2493[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_2527 = _T_2493[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_2525 = _T_2493[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_2523 = _T_2493[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2620 = {_T_2541,_T_2539,_T_2537,_T_2535,_T_2533,_T_2531,_T_2529,_T_2527,_T_2525,_T_2523}; // @[el2_lib.scala 310:69]
  wire  _T_2521 = _T_2493[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_2519 = _T_2493[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_2517 = _T_2493[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_2515 = _T_2493[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_2513 = _T_2493[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_2511 = _T_2493[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_2509 = _T_2493[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_2507 = _T_2493[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_2505 = _T_2493[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_2621 = {_T_2620,_T_2521,_T_2519,_T_2517,_T_2515,_T_2513,_T_2511,_T_2509,_T_2507,_T_2505}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_2641 = {_T_2639,_T_2630,_T_2621}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_2596 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_2602 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_2596}; // @[Cat.scala 29:58]
  wire [38:0] _T_2642 = _T_2641 ^ _T_2602; // @[el2_lib.scala 310:76]
  wire [38:0] _T_2643 = _T_2497 ? _T_2642 : _T_2602; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_2643[37:32],_T_2643[30:16],_T_2643[14:8],_T_2643[6:4],_T_2643[2]}; // @[Cat.scala 29:58]
  wire  _T_2966 = _T_2878[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_2964 = _T_2878[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_2962 = _T_2878[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_2960 = _T_2878[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_2958 = _T_2878[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_2956 = _T_2878[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_2954 = _T_2878[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_2952 = _T_2878[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_2950 = _T_2878[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_2948 = _T_2878[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3024 = {_T_2966,_T_2964,_T_2962,_T_2960,_T_2958,_T_2956,_T_2954,_T_2952,_T_2950,_T_2948}; // @[el2_lib.scala 310:69]
  wire  _T_2946 = _T_2878[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_2944 = _T_2878[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_2942 = _T_2878[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_2940 = _T_2878[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_2938 = _T_2878[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_2936 = _T_2878[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_2934 = _T_2878[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_2932 = _T_2878[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_2930 = _T_2878[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_2928 = _T_2878[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3015 = {_T_2946,_T_2944,_T_2942,_T_2940,_T_2938,_T_2936,_T_2934,_T_2932,_T_2930,_T_2928}; // @[el2_lib.scala 310:69]
  wire  _T_2926 = _T_2878[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_2924 = _T_2878[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_2922 = _T_2878[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_2920 = _T_2878[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_2918 = _T_2878[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_2916 = _T_2878[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_2914 = _T_2878[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_2912 = _T_2878[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_2910 = _T_2878[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_2908 = _T_2878[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3005 = {_T_2926,_T_2924,_T_2922,_T_2920,_T_2918,_T_2916,_T_2914,_T_2912,_T_2910,_T_2908}; // @[el2_lib.scala 310:69]
  wire  _T_2906 = _T_2878[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_2904 = _T_2878[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_2902 = _T_2878[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_2900 = _T_2878[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_2898 = _T_2878[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_2896 = _T_2878[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_2894 = _T_2878[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_2892 = _T_2878[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_2890 = _T_2878[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3006 = {_T_3005,_T_2906,_T_2904,_T_2902,_T_2900,_T_2898,_T_2896,_T_2894,_T_2892,_T_2890}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3026 = {_T_3024,_T_3015,_T_3006}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_2981 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_2987 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_2981}; // @[Cat.scala 29:58]
  wire [38:0] _T_3027 = _T_3026 ^ _T_2987; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3028 = _T_2882 ? _T_3027 : _T_2987; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3028[37:32],_T_3028[30:16],_T_3028[14:8],_T_3028[6:4],_T_3028[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 650:35]
  wire  _T_2501 = ~_T_2493[6]; // @[el2_lib.scala 303:55]
  wire  _T_2502 = _T_2495 & _T_2501; // @[el2_lib.scala 303:53]
  wire  _T_2886 = ~_T_2878[6]; // @[el2_lib.scala 303:55]
  wire  _T_2887 = _T_2880 & _T_2886; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_2502,_T_2887}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 652:53]
  wire [63:0] _T_2253 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_2254 = {iccm_dma_rdata_1_muxed,_T_2643[37:32],_T_2643[30:16],_T_2643[14:8],_T_2643[6:4],_T_2643[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 654:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 655:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 660:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 664:70]
  wire  _T_2259 = _T_1834 & _T_1823; // @[el2_ifu_mem_ctl.scala 667:65]
  wire  _T_2262 = _T_2240 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 668:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_2263 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_2265 = _T_2262 ? {{1'd0}, _T_2263} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 668:8]
  wire [31:0] _T_2266 = _T_2259 ? io_dma_mem_addr : {{16'd0}, _T_2265}; // @[el2_ifu_mem_ctl.scala 667:25]
  wire  _T_2655 = _T_2493 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_2656 = _T_2643[38] ^ _T_2655; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_2656,_T_2643[31],_T_2643[15],_T_2643[7],_T_2643[3],_T_2643[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3040 = _T_2878 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3041 = _T_3028[38] ^ _T_3040; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3041,_T_3028[31],_T_3028[15],_T_3028[7],_T_3028[3],_T_3028[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3057 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 680:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 682:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 683:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 691:62]
  wire  _T_3065 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 685:76]
  wire  _T_3066 = io_iccm_rd_ecc_single_err & _T_3065; // @[el2_ifu_mem_ctl.scala 685:74]
  wire  _T_3068 = _T_3066 & _T_317; // @[el2_ifu_mem_ctl.scala 685:104]
  wire  iccm_ecc_write_status = _T_3068 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 685:127]
  wire  _T_3069 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 686:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3069 & _T_317; // @[el2_ifu_mem_ctl.scala 686:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 690:51]
  wire [13:0] _T_3074 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 689:102]
  wire [38:0] _T_3078 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3083 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 694:41]
  wire  _T_3084 = io_ifc_fetch_req_bf & _T_3083; // @[el2_ifu_mem_ctl.scala 694:39]
  wire  _T_3085 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 694:72]
  wire  _T_3086 = _T_3084 & _T_3085; // @[el2_ifu_mem_ctl.scala 694:70]
  wire  _T_3088 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 695:34]
  wire  _T_3089 = _T_1389 & _T_3088; // @[el2_ifu_mem_ctl.scala 695:32]
  wire  _T_3092 = _T_1405 & _T_3088; // @[el2_ifu_mem_ctl.scala 696:37]
  wire  _T_3093 = _T_3089 | _T_3092; // @[el2_ifu_mem_ctl.scala 695:88]
  wire  _T_3094 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 697:19]
  wire  _T_3096 = _T_3094 & _T_3088; // @[el2_ifu_mem_ctl.scala 697:41]
  wire  _T_3097 = _T_3093 | _T_3096; // @[el2_ifu_mem_ctl.scala 696:88]
  wire  _T_3098 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 698:19]
  wire  _T_3100 = _T_3098 & _T_3088; // @[el2_ifu_mem_ctl.scala 698:35]
  wire  _T_3101 = _T_3097 | _T_3100; // @[el2_ifu_mem_ctl.scala 697:88]
  wire  _T_3104 = _T_1404 & _T_3088; // @[el2_ifu_mem_ctl.scala 699:38]
  wire  _T_3105 = _T_3101 | _T_3104; // @[el2_ifu_mem_ctl.scala 698:88]
  wire  _T_3107 = _T_1405 & miss_state_en; // @[el2_ifu_mem_ctl.scala 700:37]
  wire  _T_3108 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 700:71]
  wire  _T_3109 = _T_3107 & _T_3108; // @[el2_ifu_mem_ctl.scala 700:54]
  wire  _T_3110 = _T_3105 | _T_3109; // @[el2_ifu_mem_ctl.scala 699:57]
  wire  _T_3111 = ~_T_3110; // @[el2_ifu_mem_ctl.scala 695:5]
  wire  _T_3112 = _T_3086 & _T_3111; // @[el2_ifu_mem_ctl.scala 694:96]
  wire  _T_3113 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 701:28]
  wire  _T_3115 = _T_3113 & _T_3083; // @[el2_ifu_mem_ctl.scala 701:50]
  wire  _T_3117 = _T_3115 & _T_3085; // @[el2_ifu_mem_ctl.scala 701:81]
  wire  _T_3126 = ~_T_108; // @[el2_ifu_mem_ctl.scala 704:106]
  wire  _T_3127 = _T_1389 & _T_3126; // @[el2_ifu_mem_ctl.scala 704:104]
  wire  _T_3128 = _T_1405 | _T_3127; // @[el2_ifu_mem_ctl.scala 704:77]
  wire  _T_3132 = ~_T_51; // @[el2_ifu_mem_ctl.scala 704:172]
  wire  _T_3133 = _T_3128 & _T_3132; // @[el2_ifu_mem_ctl.scala 704:170]
  wire  _T_3134 = ~_T_3133; // @[el2_ifu_mem_ctl.scala 704:44]
  wire  _T_3138 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 707:64]
  wire  _T_3139 = ~_T_3138; // @[el2_ifu_mem_ctl.scala 707:50]
  wire  _T_3140 = _T_276 & _T_3139; // @[el2_ifu_mem_ctl.scala 707:48]
  wire  _T_3141 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 707:81]
  wire  ic_valid = _T_3140 & _T_3141; // @[el2_ifu_mem_ctl.scala 707:79]
  wire  _T_3143 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 708:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 711:14]
  wire  _T_3146 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 714:74]
  wire  _T_9288 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 788:45]
  wire  way_status_wr_en = _T_9288 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 788:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3146; // @[el2_ifu_mem_ctl.scala 714:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 716:14]
  wire [2:0] _T_3150 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 720:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 784:41]
  wire  way_status_new = _T_9288 ? replace_way_mb_any_0 : way_status_hit_new; // @[el2_ifu_mem_ctl.scala 787:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 722:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  _T_3167 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 728:93]
  wire  _T_3168 = _T_3167 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:102]
  wire  _T_3169 = _T_3168 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3171 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 728:93]
  wire  _T_3172 = _T_3171 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:102]
  wire  _T_3173 = _T_3172 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3175 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 728:93]
  wire  _T_3176 = _T_3175 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:102]
  wire  _T_3177 = _T_3176 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3179 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 728:93]
  wire  _T_3180 = _T_3179 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:102]
  wire  _T_3181 = _T_3180 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3183 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 728:93]
  wire  _T_3184 = _T_3183 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:102]
  wire  _T_3185 = _T_3184 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3187 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 728:93]
  wire  _T_3188 = _T_3187 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:102]
  wire  _T_3189 = _T_3188 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3191 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 728:93]
  wire  _T_3192 = _T_3191 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:102]
  wire  _T_3193 = _T_3192 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3195 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 728:93]
  wire  _T_3196 = _T_3195 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:102]
  wire  _T_3197 = _T_3196 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3201 = _T_3168 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3205 = _T_3172 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3209 = _T_3176 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3213 = _T_3180 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3217 = _T_3184 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3221 = _T_3188 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3225 = _T_3192 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3229 = _T_3196 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3233 = _T_3168 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3237 = _T_3172 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3241 = _T_3176 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3245 = _T_3180 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3249 = _T_3184 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3253 = _T_3188 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3257 = _T_3192 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3261 = _T_3196 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3265 = _T_3168 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3269 = _T_3172 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3273 = _T_3176 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3277 = _T_3180 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3281 = _T_3184 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3285 = _T_3188 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3289 = _T_3192 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3293 = _T_3196 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3297 = _T_3168 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3301 = _T_3172 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3305 = _T_3176 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3309 = _T_3180 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3313 = _T_3184 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3317 = _T_3188 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3321 = _T_3192 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3325 = _T_3196 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3329 = _T_3168 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3333 = _T_3172 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3337 = _T_3176 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3341 = _T_3180 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3345 = _T_3184 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3349 = _T_3188 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3353 = _T_3192 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3357 = _T_3196 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3361 = _T_3168 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3365 = _T_3172 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3369 = _T_3176 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3373 = _T_3180 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3377 = _T_3184 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3381 = _T_3188 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3385 = _T_3192 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3389 = _T_3196 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3393 = _T_3168 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3397 = _T_3172 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3401 = _T_3176 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3405 = _T_3180 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3409 = _T_3184 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3413 = _T_3188 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3417 = _T_3192 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3421 = _T_3196 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3425 = _T_3168 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3429 = _T_3172 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3433 = _T_3176 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3437 = _T_3180 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3441 = _T_3184 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3445 = _T_3188 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3449 = _T_3192 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3453 = _T_3196 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3457 = _T_3168 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3461 = _T_3172 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3465 = _T_3176 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3469 = _T_3180 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3473 = _T_3184 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3477 = _T_3188 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3481 = _T_3192 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3485 = _T_3196 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3489 = _T_3168 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3493 = _T_3172 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3497 = _T_3176 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3501 = _T_3180 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3505 = _T_3184 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3509 = _T_3188 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3513 = _T_3192 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3517 = _T_3196 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3521 = _T_3168 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3525 = _T_3172 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3529 = _T_3176 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3533 = _T_3180 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3537 = _T_3184 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3541 = _T_3188 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3545 = _T_3192 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3549 = _T_3196 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3553 = _T_3168 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3557 = _T_3172 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3561 = _T_3176 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3565 = _T_3180 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3569 = _T_3184 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3573 = _T_3188 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3577 = _T_3192 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3581 = _T_3196 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3585 = _T_3168 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3589 = _T_3172 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3593 = _T_3176 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3597 = _T_3180 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3601 = _T_3184 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3605 = _T_3188 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3609 = _T_3192 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3613 = _T_3196 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3617 = _T_3168 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3621 = _T_3172 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3625 = _T_3176 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3629 = _T_3180 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3633 = _T_3184 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3637 = _T_3188 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3641 = _T_3192 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3645 = _T_3196 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3649 = _T_3168 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3653 = _T_3172 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3657 = _T_3176 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3661 = _T_3180 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3665 = _T_3184 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3669 = _T_3188 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3673 = _T_3192 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_3677 = _T_3196 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:124]
  wire  _T_9294 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 791:84]
  wire  _T_9295 = _T_9294 & miss_pending; // @[el2_ifu_mem_ctl.scala 791:108]
  wire  bus_wren_last_1 = _T_9295 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 791:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 792:84]
  wire  _T_9297 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 793:73]
  wire  _T_9292 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 791:84]
  wire  _T_9293 = _T_9292 & miss_pending; // @[el2_ifu_mem_ctl.scala 791:108]
  wire  bus_wren_last_0 = _T_9293 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 791:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 792:84]
  wire  _T_9296 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 793:73]
  wire [1:0] ifu_tag_wren = {_T_9297,_T_9296}; // @[Cat.scala 29:58]
  wire [1:0] _T_9331 = _T_3146 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9331 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 826:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 737:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 739:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 743:14]
  wire  _T_4326 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 747:82]
  wire  _T_4328 = _T_4326 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 747:91]
  wire  _T_4330 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 748:74]
  wire  _T_4332 = _T_4330 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 748:83]
  wire  _T_4333 = _T_4328 | _T_4332; // @[el2_ifu_mem_ctl.scala 747:113]
  wire  _T_4334 = _T_4333 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:106]
  wire  _T_4338 = _T_4326 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 747:91]
  wire  _T_4342 = _T_4330 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 748:83]
  wire  _T_4343 = _T_4338 | _T_4342; // @[el2_ifu_mem_ctl.scala 747:113]
  wire  _T_4344 = _T_4343 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:106]
  wire [1:0] tag_valid_clken_0 = {_T_4334,_T_4344}; // @[Cat.scala 29:58]
  wire  _T_4346 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 747:82]
  wire  _T_4348 = _T_4346 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 747:91]
  wire  _T_4350 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 748:74]
  wire  _T_4352 = _T_4350 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 748:83]
  wire  _T_4353 = _T_4348 | _T_4352; // @[el2_ifu_mem_ctl.scala 747:113]
  wire  _T_4354 = _T_4353 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:106]
  wire  _T_4358 = _T_4346 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 747:91]
  wire  _T_4362 = _T_4350 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 748:83]
  wire  _T_4363 = _T_4358 | _T_4362; // @[el2_ifu_mem_ctl.scala 747:113]
  wire  _T_4364 = _T_4363 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:106]
  wire [1:0] tag_valid_clken_1 = {_T_4354,_T_4364}; // @[Cat.scala 29:58]
  wire  _T_4366 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 747:82]
  wire  _T_4368 = _T_4366 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 747:91]
  wire  _T_4370 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 748:74]
  wire  _T_4372 = _T_4370 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 748:83]
  wire  _T_4373 = _T_4368 | _T_4372; // @[el2_ifu_mem_ctl.scala 747:113]
  wire  _T_4374 = _T_4373 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:106]
  wire  _T_4378 = _T_4366 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 747:91]
  wire  _T_4382 = _T_4370 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 748:83]
  wire  _T_4383 = _T_4378 | _T_4382; // @[el2_ifu_mem_ctl.scala 747:113]
  wire  _T_4384 = _T_4383 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:106]
  wire [1:0] tag_valid_clken_2 = {_T_4374,_T_4384}; // @[Cat.scala 29:58]
  wire  _T_4386 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 747:82]
  wire  _T_4388 = _T_4386 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 747:91]
  wire  _T_4390 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 748:74]
  wire  _T_4392 = _T_4390 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 748:83]
  wire  _T_4393 = _T_4388 | _T_4392; // @[el2_ifu_mem_ctl.scala 747:113]
  wire  _T_4394 = _T_4393 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:106]
  wire  _T_4398 = _T_4386 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 747:91]
  wire  _T_4402 = _T_4390 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 748:83]
  wire  _T_4403 = _T_4398 | _T_4402; // @[el2_ifu_mem_ctl.scala 747:113]
  wire  _T_4404 = _T_4403 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:106]
  wire [1:0] tag_valid_clken_3 = {_T_4394,_T_4404}; // @[Cat.scala 29:58]
  wire  _T_4407 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 753:64]
  wire  _T_4408 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 753:91]
  wire  _T_4409 = _T_4407 & _T_4408; // @[el2_ifu_mem_ctl.scala 753:89]
  wire  _T_4412 = _T_3679 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4413 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4415 = _T_4413 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4417 = _T_4415 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4418 = _T_4412 | _T_4417; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4428 = _T_3683 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4429 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4431 = _T_4429 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4433 = _T_4431 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4434 = _T_4428 | _T_4433; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4444 = _T_3687 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4445 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4447 = _T_4445 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4449 = _T_4447 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4450 = _T_4444 | _T_4449; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4460 = _T_3691 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4461 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4463 = _T_4461 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4465 = _T_4463 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4466 = _T_4460 | _T_4465; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4476 = _T_3695 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4477 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4479 = _T_4477 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4481 = _T_4479 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4482 = _T_4476 | _T_4481; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4492 = _T_3699 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4493 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4495 = _T_4493 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4497 = _T_4495 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4498 = _T_4492 | _T_4497; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4508 = _T_3703 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4509 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4511 = _T_4509 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4513 = _T_4511 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4514 = _T_4508 | _T_4513; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4524 = _T_3707 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4525 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4527 = _T_4525 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4529 = _T_4527 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4530 = _T_4524 | _T_4529; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4540 = _T_3711 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4541 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4543 = _T_4541 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4545 = _T_4543 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4546 = _T_4540 | _T_4545; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4556 = _T_3715 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4557 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4559 = _T_4557 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4561 = _T_4559 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4562 = _T_4556 | _T_4561; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4572 = _T_3719 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4573 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4575 = _T_4573 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4577 = _T_4575 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4578 = _T_4572 | _T_4577; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4588 = _T_3723 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4589 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4591 = _T_4589 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4593 = _T_4591 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4594 = _T_4588 | _T_4593; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4604 = _T_3727 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4605 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4607 = _T_4605 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4609 = _T_4607 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4610 = _T_4604 | _T_4609; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4620 = _T_3731 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4621 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4623 = _T_4621 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4625 = _T_4623 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4626 = _T_4620 | _T_4625; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4636 = _T_3735 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4637 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4639 = _T_4637 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4641 = _T_4639 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4642 = _T_4636 | _T_4641; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4652 = _T_3739 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4653 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4655 = _T_4653 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4657 = _T_4655 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4658 = _T_4652 | _T_4657; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4668 = _T_3743 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4669 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4671 = _T_4669 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4673 = _T_4671 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4674 = _T_4668 | _T_4673; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4684 = _T_3747 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4685 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4687 = _T_4685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4689 = _T_4687 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4690 = _T_4684 | _T_4689; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4700 = _T_3751 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4701 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4703 = _T_4701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4705 = _T_4703 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4706 = _T_4700 | _T_4705; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4716 = _T_3755 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4717 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4719 = _T_4717 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4721 = _T_4719 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4722 = _T_4716 | _T_4721; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4732 = _T_3759 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4733 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4735 = _T_4733 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4737 = _T_4735 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4738 = _T_4732 | _T_4737; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4748 = _T_3763 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4749 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4751 = _T_4749 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4753 = _T_4751 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4754 = _T_4748 | _T_4753; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4764 = _T_3767 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4765 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4767 = _T_4765 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4769 = _T_4767 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4770 = _T_4764 | _T_4769; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4780 = _T_3771 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4781 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4783 = _T_4781 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4785 = _T_4783 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4786 = _T_4780 | _T_4785; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4796 = _T_3775 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4797 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4799 = _T_4797 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4801 = _T_4799 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4802 = _T_4796 | _T_4801; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4812 = _T_3779 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4813 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4815 = _T_4813 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4817 = _T_4815 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4818 = _T_4812 | _T_4817; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4828 = _T_3783 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4829 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4831 = _T_4829 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4833 = _T_4831 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4834 = _T_4828 | _T_4833; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4844 = _T_3787 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4845 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4847 = _T_4845 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4849 = _T_4847 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4850 = _T_4844 | _T_4849; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4860 = _T_3791 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4861 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4863 = _T_4861 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4865 = _T_4863 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4866 = _T_4860 | _T_4865; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4876 = _T_3795 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4877 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4879 = _T_4877 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4881 = _T_4879 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4882 = _T_4876 | _T_4881; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4892 = _T_3799 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4893 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4895 = _T_4893 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4897 = _T_4895 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4898 = _T_4892 | _T_4897; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4908 = _T_3803 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4909 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_4911 = _T_4909 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4913 = _T_4911 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4914 = _T_4908 | _T_4913; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4924 = _T_3679 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4927 = _T_4413 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4929 = _T_4927 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4930 = _T_4924 | _T_4929; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4940 = _T_3683 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4943 = _T_4429 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4945 = _T_4943 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4946 = _T_4940 | _T_4945; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4956 = _T_3687 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4959 = _T_4445 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4961 = _T_4959 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4962 = _T_4956 | _T_4961; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4972 = _T_3691 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4975 = _T_4461 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4977 = _T_4975 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4978 = _T_4972 | _T_4977; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_4988 = _T_3695 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_4991 = _T_4477 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_4993 = _T_4991 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_4994 = _T_4988 | _T_4993; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5004 = _T_3699 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5007 = _T_4493 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5009 = _T_5007 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5010 = _T_5004 | _T_5009; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5020 = _T_3703 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5023 = _T_4509 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5025 = _T_5023 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5026 = _T_5020 | _T_5025; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5036 = _T_3707 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5039 = _T_4525 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5041 = _T_5039 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5042 = _T_5036 | _T_5041; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5052 = _T_3711 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5055 = _T_4541 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5057 = _T_5055 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5058 = _T_5052 | _T_5057; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5068 = _T_3715 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5071 = _T_4557 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5073 = _T_5071 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5074 = _T_5068 | _T_5073; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5084 = _T_3719 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5087 = _T_4573 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5089 = _T_5087 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5090 = _T_5084 | _T_5089; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5100 = _T_3723 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5103 = _T_4589 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5105 = _T_5103 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5106 = _T_5100 | _T_5105; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5116 = _T_3727 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5119 = _T_4605 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5121 = _T_5119 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5122 = _T_5116 | _T_5121; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5132 = _T_3731 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5135 = _T_4621 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5137 = _T_5135 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5138 = _T_5132 | _T_5137; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5148 = _T_3735 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5151 = _T_4637 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5153 = _T_5151 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5154 = _T_5148 | _T_5153; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5164 = _T_3739 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5167 = _T_4653 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5169 = _T_5167 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5170 = _T_5164 | _T_5169; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5180 = _T_3743 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5183 = _T_4669 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5185 = _T_5183 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5186 = _T_5180 | _T_5185; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5196 = _T_3747 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5199 = _T_4685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5201 = _T_5199 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5202 = _T_5196 | _T_5201; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5212 = _T_3751 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5215 = _T_4701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5217 = _T_5215 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5218 = _T_5212 | _T_5217; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5228 = _T_3755 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5231 = _T_4717 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5233 = _T_5231 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5234 = _T_5228 | _T_5233; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5244 = _T_3759 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5247 = _T_4733 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5249 = _T_5247 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5250 = _T_5244 | _T_5249; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5260 = _T_3763 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5263 = _T_4749 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5265 = _T_5263 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5266 = _T_5260 | _T_5265; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5276 = _T_3767 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5279 = _T_4765 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5281 = _T_5279 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5282 = _T_5276 | _T_5281; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5292 = _T_3771 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5295 = _T_4781 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5297 = _T_5295 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5298 = _T_5292 | _T_5297; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5308 = _T_3775 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5311 = _T_4797 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5313 = _T_5311 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5314 = _T_5308 | _T_5313; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5324 = _T_3779 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5327 = _T_4813 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5329 = _T_5327 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5330 = _T_5324 | _T_5329; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5340 = _T_3783 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5343 = _T_4829 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5345 = _T_5343 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5346 = _T_5340 | _T_5345; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5356 = _T_3787 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5359 = _T_4845 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5361 = _T_5359 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5362 = _T_5356 | _T_5361; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5372 = _T_3791 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5375 = _T_4861 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5377 = _T_5375 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5378 = _T_5372 | _T_5377; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5388 = _T_3795 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5391 = _T_4877 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5393 = _T_5391 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5394 = _T_5388 | _T_5393; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5404 = _T_3799 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5407 = _T_4893 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5409 = _T_5407 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5410 = _T_5404 | _T_5409; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5420 = _T_3803 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5423 = _T_4909 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5425 = _T_5423 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5426 = _T_5420 | _T_5425; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5436 = _T_3807 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5437 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5439 = _T_5437 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5441 = _T_5439 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5442 = _T_5436 | _T_5441; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5452 = _T_3811 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5453 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5455 = _T_5453 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5457 = _T_5455 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5458 = _T_5452 | _T_5457; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5468 = _T_3815 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5469 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5471 = _T_5469 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5473 = _T_5471 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5474 = _T_5468 | _T_5473; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5484 = _T_3819 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5485 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5487 = _T_5485 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5489 = _T_5487 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5490 = _T_5484 | _T_5489; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5500 = _T_3823 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5501 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5503 = _T_5501 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5505 = _T_5503 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5506 = _T_5500 | _T_5505; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5516 = _T_3827 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5517 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5519 = _T_5517 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5521 = _T_5519 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5522 = _T_5516 | _T_5521; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5532 = _T_3831 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5533 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5535 = _T_5533 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5537 = _T_5535 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5538 = _T_5532 | _T_5537; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5548 = _T_3835 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5549 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5551 = _T_5549 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5553 = _T_5551 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5554 = _T_5548 | _T_5553; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5564 = _T_3839 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5565 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5567 = _T_5565 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5569 = _T_5567 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5570 = _T_5564 | _T_5569; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5580 = _T_3843 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5581 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5583 = _T_5581 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5585 = _T_5583 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5586 = _T_5580 | _T_5585; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5596 = _T_3847 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5597 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5599 = _T_5597 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5601 = _T_5599 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5602 = _T_5596 | _T_5601; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5612 = _T_3851 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5613 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5615 = _T_5613 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5617 = _T_5615 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5618 = _T_5612 | _T_5617; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5628 = _T_3855 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5629 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5631 = _T_5629 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5633 = _T_5631 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5634 = _T_5628 | _T_5633; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5644 = _T_3859 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5645 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5647 = _T_5645 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5649 = _T_5647 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5650 = _T_5644 | _T_5649; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5660 = _T_3863 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5661 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5663 = _T_5661 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5665 = _T_5663 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5666 = _T_5660 | _T_5665; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5676 = _T_3867 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5677 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5679 = _T_5677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5681 = _T_5679 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5682 = _T_5676 | _T_5681; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5692 = _T_3871 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5693 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5695 = _T_5693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5697 = _T_5695 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5698 = _T_5692 | _T_5697; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5708 = _T_3875 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5709 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5711 = _T_5709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5713 = _T_5711 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5714 = _T_5708 | _T_5713; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5724 = _T_3879 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5725 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5727 = _T_5725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5729 = _T_5727 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5730 = _T_5724 | _T_5729; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5740 = _T_3883 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5741 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5743 = _T_5741 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5745 = _T_5743 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5746 = _T_5740 | _T_5745; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5756 = _T_3887 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5757 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5759 = _T_5757 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5761 = _T_5759 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5762 = _T_5756 | _T_5761; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5772 = _T_3891 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5773 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5775 = _T_5773 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5777 = _T_5775 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5778 = _T_5772 | _T_5777; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5788 = _T_3895 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5789 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5791 = _T_5789 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5793 = _T_5791 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5794 = _T_5788 | _T_5793; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5804 = _T_3899 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5805 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5807 = _T_5805 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5809 = _T_5807 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5810 = _T_5804 | _T_5809; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5820 = _T_3903 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5821 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5823 = _T_5821 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5825 = _T_5823 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5826 = _T_5820 | _T_5825; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5836 = _T_3907 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5837 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5839 = _T_5837 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5841 = _T_5839 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5842 = _T_5836 | _T_5841; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5852 = _T_3911 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5853 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5855 = _T_5853 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5857 = _T_5855 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5858 = _T_5852 | _T_5857; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5868 = _T_3915 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5869 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5871 = _T_5869 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5873 = _T_5871 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5874 = _T_5868 | _T_5873; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5884 = _T_3919 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5885 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5887 = _T_5885 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5889 = _T_5887 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5890 = _T_5884 | _T_5889; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5900 = _T_3923 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5901 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5903 = _T_5901 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5905 = _T_5903 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5906 = _T_5900 | _T_5905; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5916 = _T_3927 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5917 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5919 = _T_5917 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5921 = _T_5919 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5922 = _T_5916 | _T_5921; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5932 = _T_3931 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5933 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_5935 = _T_5933 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5937 = _T_5935 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5938 = _T_5932 | _T_5937; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5948 = _T_3807 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5951 = _T_5437 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5953 = _T_5951 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5954 = _T_5948 | _T_5953; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5964 = _T_3811 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5967 = _T_5453 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5969 = _T_5967 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5970 = _T_5964 | _T_5969; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5980 = _T_3815 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5983 = _T_5469 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_5985 = _T_5983 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_5986 = _T_5980 | _T_5985; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_5996 = _T_3819 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_5999 = _T_5485 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6001 = _T_5999 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6002 = _T_5996 | _T_6001; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6012 = _T_3823 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6015 = _T_5501 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6017 = _T_6015 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6018 = _T_6012 | _T_6017; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6028 = _T_3827 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6031 = _T_5517 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6033 = _T_6031 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6034 = _T_6028 | _T_6033; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6044 = _T_3831 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6047 = _T_5533 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6049 = _T_6047 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6050 = _T_6044 | _T_6049; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6060 = _T_3835 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6063 = _T_5549 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6065 = _T_6063 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6066 = _T_6060 | _T_6065; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6076 = _T_3839 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6079 = _T_5565 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6081 = _T_6079 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6082 = _T_6076 | _T_6081; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6092 = _T_3843 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6095 = _T_5581 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6097 = _T_6095 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6098 = _T_6092 | _T_6097; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6108 = _T_3847 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6111 = _T_5597 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6113 = _T_6111 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6114 = _T_6108 | _T_6113; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6124 = _T_3851 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6127 = _T_5613 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6129 = _T_6127 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6130 = _T_6124 | _T_6129; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6140 = _T_3855 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6143 = _T_5629 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6145 = _T_6143 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6146 = _T_6140 | _T_6145; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6156 = _T_3859 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6159 = _T_5645 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6161 = _T_6159 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6162 = _T_6156 | _T_6161; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6172 = _T_3863 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6175 = _T_5661 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6177 = _T_6175 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6178 = _T_6172 | _T_6177; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6188 = _T_3867 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6191 = _T_5677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6193 = _T_6191 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6194 = _T_6188 | _T_6193; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6204 = _T_3871 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6207 = _T_5693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6209 = _T_6207 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6210 = _T_6204 | _T_6209; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6220 = _T_3875 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6223 = _T_5709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6225 = _T_6223 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6226 = _T_6220 | _T_6225; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6236 = _T_3879 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6239 = _T_5725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6241 = _T_6239 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6242 = _T_6236 | _T_6241; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6252 = _T_3883 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6255 = _T_5741 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6257 = _T_6255 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6258 = _T_6252 | _T_6257; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6268 = _T_3887 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6271 = _T_5757 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6273 = _T_6271 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6274 = _T_6268 | _T_6273; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6284 = _T_3891 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6287 = _T_5773 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6289 = _T_6287 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6290 = _T_6284 | _T_6289; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6300 = _T_3895 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6303 = _T_5789 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6305 = _T_6303 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6306 = _T_6300 | _T_6305; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6316 = _T_3899 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6319 = _T_5805 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6321 = _T_6319 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6322 = _T_6316 | _T_6321; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6332 = _T_3903 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6335 = _T_5821 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6337 = _T_6335 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6338 = _T_6332 | _T_6337; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6348 = _T_3907 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6351 = _T_5837 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6353 = _T_6351 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6354 = _T_6348 | _T_6353; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6364 = _T_3911 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6367 = _T_5853 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6369 = _T_6367 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6370 = _T_6364 | _T_6369; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6380 = _T_3915 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6383 = _T_5869 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6385 = _T_6383 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6386 = _T_6380 | _T_6385; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6396 = _T_3919 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6399 = _T_5885 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6401 = _T_6399 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6402 = _T_6396 | _T_6401; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6412 = _T_3923 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6415 = _T_5901 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6417 = _T_6415 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6418 = _T_6412 | _T_6417; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6428 = _T_3927 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6431 = _T_5917 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6433 = _T_6431 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6434 = _T_6428 | _T_6433; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6444 = _T_3931 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6447 = _T_5933 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6449 = _T_6447 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6450 = _T_6444 | _T_6449; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6460 = _T_3935 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire [6:0] _GEN_797 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6461 = _GEN_797 == 7'h40; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6463 = _T_6461 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6465 = _T_6463 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6466 = _T_6460 | _T_6465; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6476 = _T_3939 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6477 = _GEN_797 == 7'h41; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6479 = _T_6477 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6481 = _T_6479 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6482 = _T_6476 | _T_6481; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6492 = _T_3943 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6493 = _GEN_797 == 7'h42; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6495 = _T_6493 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6497 = _T_6495 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6498 = _T_6492 | _T_6497; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6508 = _T_3947 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6509 = _GEN_797 == 7'h43; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6511 = _T_6509 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6513 = _T_6511 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6514 = _T_6508 | _T_6513; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6524 = _T_3951 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6525 = _GEN_797 == 7'h44; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6527 = _T_6525 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6529 = _T_6527 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6530 = _T_6524 | _T_6529; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6540 = _T_3955 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6541 = _GEN_797 == 7'h45; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6543 = _T_6541 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6545 = _T_6543 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6546 = _T_6540 | _T_6545; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6556 = _T_3959 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6557 = _GEN_797 == 7'h46; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6559 = _T_6557 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6561 = _T_6559 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6562 = _T_6556 | _T_6561; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6572 = _T_3963 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6573 = _GEN_797 == 7'h47; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6575 = _T_6573 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6577 = _T_6575 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6578 = _T_6572 | _T_6577; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6588 = _T_3967 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6589 = _GEN_797 == 7'h48; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6591 = _T_6589 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6593 = _T_6591 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6594 = _T_6588 | _T_6593; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6604 = _T_3971 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6605 = _GEN_797 == 7'h49; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6607 = _T_6605 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6609 = _T_6607 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6610 = _T_6604 | _T_6609; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6620 = _T_3975 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6621 = _GEN_797 == 7'h4a; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6623 = _T_6621 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6625 = _T_6623 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6626 = _T_6620 | _T_6625; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6636 = _T_3979 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6637 = _GEN_797 == 7'h4b; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6639 = _T_6637 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6641 = _T_6639 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6642 = _T_6636 | _T_6641; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6652 = _T_3983 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6653 = _GEN_797 == 7'h4c; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6655 = _T_6653 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6657 = _T_6655 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6658 = _T_6652 | _T_6657; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6668 = _T_3987 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6669 = _GEN_797 == 7'h4d; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6671 = _T_6669 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6673 = _T_6671 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6674 = _T_6668 | _T_6673; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6684 = _T_3991 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6685 = _GEN_797 == 7'h4e; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6687 = _T_6685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6689 = _T_6687 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6690 = _T_6684 | _T_6689; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6700 = _T_3995 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6701 = _GEN_797 == 7'h4f; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6703 = _T_6701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6705 = _T_6703 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6706 = _T_6700 | _T_6705; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6716 = _T_3999 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6717 = _GEN_797 == 7'h50; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6719 = _T_6717 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6721 = _T_6719 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6722 = _T_6716 | _T_6721; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6732 = _T_4003 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6733 = _GEN_797 == 7'h51; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6735 = _T_6733 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6737 = _T_6735 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6738 = _T_6732 | _T_6737; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6748 = _T_4007 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6749 = _GEN_797 == 7'h52; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6751 = _T_6749 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6753 = _T_6751 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6754 = _T_6748 | _T_6753; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6764 = _T_4011 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6765 = _GEN_797 == 7'h53; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6767 = _T_6765 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6769 = _T_6767 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6770 = _T_6764 | _T_6769; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6780 = _T_4015 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6781 = _GEN_797 == 7'h54; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6783 = _T_6781 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6785 = _T_6783 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6786 = _T_6780 | _T_6785; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6796 = _T_4019 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6797 = _GEN_797 == 7'h55; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6799 = _T_6797 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6801 = _T_6799 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6802 = _T_6796 | _T_6801; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6812 = _T_4023 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6813 = _GEN_797 == 7'h56; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6815 = _T_6813 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6817 = _T_6815 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6818 = _T_6812 | _T_6817; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6828 = _T_4027 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6829 = _GEN_797 == 7'h57; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6831 = _T_6829 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6833 = _T_6831 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6834 = _T_6828 | _T_6833; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6844 = _T_4031 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6845 = _GEN_797 == 7'h58; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6847 = _T_6845 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6849 = _T_6847 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6850 = _T_6844 | _T_6849; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6860 = _T_4035 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6861 = _GEN_797 == 7'h59; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6863 = _T_6861 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6865 = _T_6863 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6866 = _T_6860 | _T_6865; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6876 = _T_4039 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6877 = _GEN_797 == 7'h5a; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6879 = _T_6877 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6881 = _T_6879 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6882 = _T_6876 | _T_6881; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6892 = _T_4043 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6893 = _GEN_797 == 7'h5b; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6895 = _T_6893 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6897 = _T_6895 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6898 = _T_6892 | _T_6897; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6908 = _T_4047 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6909 = _GEN_797 == 7'h5c; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6911 = _T_6909 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6913 = _T_6911 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6914 = _T_6908 | _T_6913; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6924 = _T_4051 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6925 = _GEN_797 == 7'h5d; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6927 = _T_6925 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6929 = _T_6927 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6930 = _T_6924 | _T_6929; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6940 = _T_4055 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6941 = _GEN_797 == 7'h5e; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6943 = _T_6941 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6945 = _T_6943 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6946 = _T_6940 | _T_6945; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6956 = _T_4059 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6957 = _GEN_797 == 7'h5f; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_6959 = _T_6957 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6961 = _T_6959 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6962 = _T_6956 | _T_6961; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6972 = _T_3935 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6975 = _T_6461 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6977 = _T_6975 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6978 = _T_6972 | _T_6977; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_6988 = _T_3939 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_6991 = _T_6477 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_6993 = _T_6991 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_6994 = _T_6988 | _T_6993; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7004 = _T_3943 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7007 = _T_6493 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7009 = _T_7007 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7010 = _T_7004 | _T_7009; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7020 = _T_3947 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7023 = _T_6509 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7025 = _T_7023 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7026 = _T_7020 | _T_7025; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7036 = _T_3951 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7039 = _T_6525 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7041 = _T_7039 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7042 = _T_7036 | _T_7041; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7052 = _T_3955 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7055 = _T_6541 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7057 = _T_7055 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7058 = _T_7052 | _T_7057; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7068 = _T_3959 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7071 = _T_6557 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7073 = _T_7071 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7074 = _T_7068 | _T_7073; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7084 = _T_3963 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7087 = _T_6573 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7089 = _T_7087 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7090 = _T_7084 | _T_7089; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7100 = _T_3967 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7103 = _T_6589 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7105 = _T_7103 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7106 = _T_7100 | _T_7105; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7116 = _T_3971 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7119 = _T_6605 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7121 = _T_7119 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7122 = _T_7116 | _T_7121; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7132 = _T_3975 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7135 = _T_6621 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7137 = _T_7135 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7138 = _T_7132 | _T_7137; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7148 = _T_3979 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7151 = _T_6637 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7153 = _T_7151 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7154 = _T_7148 | _T_7153; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7164 = _T_3983 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7167 = _T_6653 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7169 = _T_7167 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7170 = _T_7164 | _T_7169; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7180 = _T_3987 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7183 = _T_6669 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7185 = _T_7183 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7186 = _T_7180 | _T_7185; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7196 = _T_3991 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7199 = _T_6685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7201 = _T_7199 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7202 = _T_7196 | _T_7201; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7212 = _T_3995 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7215 = _T_6701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7217 = _T_7215 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7218 = _T_7212 | _T_7217; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7228 = _T_3999 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7231 = _T_6717 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7233 = _T_7231 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7234 = _T_7228 | _T_7233; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7244 = _T_4003 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7247 = _T_6733 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7249 = _T_7247 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7250 = _T_7244 | _T_7249; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7260 = _T_4007 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7263 = _T_6749 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7265 = _T_7263 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7266 = _T_7260 | _T_7265; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7276 = _T_4011 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7279 = _T_6765 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7281 = _T_7279 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7282 = _T_7276 | _T_7281; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7292 = _T_4015 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7295 = _T_6781 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7297 = _T_7295 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7298 = _T_7292 | _T_7297; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7308 = _T_4019 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7311 = _T_6797 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7313 = _T_7311 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7314 = _T_7308 | _T_7313; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7324 = _T_4023 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7327 = _T_6813 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7329 = _T_7327 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7330 = _T_7324 | _T_7329; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7340 = _T_4027 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7343 = _T_6829 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7345 = _T_7343 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7346 = _T_7340 | _T_7345; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7356 = _T_4031 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7359 = _T_6845 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7361 = _T_7359 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7362 = _T_7356 | _T_7361; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7372 = _T_4035 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7375 = _T_6861 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7377 = _T_7375 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7378 = _T_7372 | _T_7377; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7388 = _T_4039 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7391 = _T_6877 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7393 = _T_7391 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7394 = _T_7388 | _T_7393; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7404 = _T_4043 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7407 = _T_6893 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7409 = _T_7407 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7410 = _T_7404 | _T_7409; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7420 = _T_4047 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7423 = _T_6909 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7425 = _T_7423 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7426 = _T_7420 | _T_7425; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7436 = _T_4051 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7439 = _T_6925 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7441 = _T_7439 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7442 = _T_7436 | _T_7441; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7452 = _T_4055 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7455 = _T_6941 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7457 = _T_7455 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7458 = _T_7452 | _T_7457; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7468 = _T_4059 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7471 = _T_6957 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7473 = _T_7471 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7474 = _T_7468 | _T_7473; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7484 = _T_4063 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7485 = _GEN_797 == 7'h60; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7487 = _T_7485 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7489 = _T_7487 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7490 = _T_7484 | _T_7489; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7500 = _T_4067 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7501 = _GEN_797 == 7'h61; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7503 = _T_7501 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7505 = _T_7503 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7506 = _T_7500 | _T_7505; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7516 = _T_4071 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7517 = _GEN_797 == 7'h62; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7519 = _T_7517 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7521 = _T_7519 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7522 = _T_7516 | _T_7521; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7532 = _T_4075 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7533 = _GEN_797 == 7'h63; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7535 = _T_7533 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7537 = _T_7535 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7538 = _T_7532 | _T_7537; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7548 = _T_4079 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7549 = _GEN_797 == 7'h64; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7551 = _T_7549 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7553 = _T_7551 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7554 = _T_7548 | _T_7553; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7564 = _T_4083 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7565 = _GEN_797 == 7'h65; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7567 = _T_7565 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7569 = _T_7567 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7570 = _T_7564 | _T_7569; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7580 = _T_4087 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7581 = _GEN_797 == 7'h66; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7583 = _T_7581 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7585 = _T_7583 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7586 = _T_7580 | _T_7585; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7596 = _T_4091 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7597 = _GEN_797 == 7'h67; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7599 = _T_7597 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7601 = _T_7599 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7602 = _T_7596 | _T_7601; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7612 = _T_4095 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7613 = _GEN_797 == 7'h68; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7615 = _T_7613 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7617 = _T_7615 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7618 = _T_7612 | _T_7617; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7628 = _T_4099 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7629 = _GEN_797 == 7'h69; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7631 = _T_7629 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7633 = _T_7631 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7634 = _T_7628 | _T_7633; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7644 = _T_4103 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7645 = _GEN_797 == 7'h6a; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7647 = _T_7645 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7649 = _T_7647 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7650 = _T_7644 | _T_7649; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7660 = _T_4107 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7661 = _GEN_797 == 7'h6b; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7663 = _T_7661 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7665 = _T_7663 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7666 = _T_7660 | _T_7665; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7676 = _T_4111 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7677 = _GEN_797 == 7'h6c; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7679 = _T_7677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7681 = _T_7679 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7682 = _T_7676 | _T_7681; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7692 = _T_4115 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7693 = _GEN_797 == 7'h6d; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7695 = _T_7693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7697 = _T_7695 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7698 = _T_7692 | _T_7697; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7708 = _T_4119 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7709 = _GEN_797 == 7'h6e; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7711 = _T_7709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7713 = _T_7711 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7714 = _T_7708 | _T_7713; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7724 = _T_4123 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7725 = _GEN_797 == 7'h6f; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7727 = _T_7725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7729 = _T_7727 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7730 = _T_7724 | _T_7729; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7740 = _T_4127 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7741 = _GEN_797 == 7'h70; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7743 = _T_7741 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7745 = _T_7743 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7746 = _T_7740 | _T_7745; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7756 = _T_4131 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7757 = _GEN_797 == 7'h71; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7759 = _T_7757 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7761 = _T_7759 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7762 = _T_7756 | _T_7761; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7772 = _T_4135 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7773 = _GEN_797 == 7'h72; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7775 = _T_7773 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7777 = _T_7775 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7778 = _T_7772 | _T_7777; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7788 = _T_4139 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7789 = _GEN_797 == 7'h73; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7791 = _T_7789 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7793 = _T_7791 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7794 = _T_7788 | _T_7793; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7804 = _T_4143 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7805 = _GEN_797 == 7'h74; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7807 = _T_7805 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7809 = _T_7807 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7810 = _T_7804 | _T_7809; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7820 = _T_4147 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7821 = _GEN_797 == 7'h75; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7823 = _T_7821 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7825 = _T_7823 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7826 = _T_7820 | _T_7825; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7836 = _T_4151 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7837 = _GEN_797 == 7'h76; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7839 = _T_7837 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7841 = _T_7839 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7842 = _T_7836 | _T_7841; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7852 = _T_4155 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7853 = _GEN_797 == 7'h77; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7855 = _T_7853 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7857 = _T_7855 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7858 = _T_7852 | _T_7857; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7868 = _T_4159 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7869 = _GEN_797 == 7'h78; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7871 = _T_7869 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7873 = _T_7871 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7874 = _T_7868 | _T_7873; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7884 = _T_4163 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7885 = _GEN_797 == 7'h79; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7887 = _T_7885 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7889 = _T_7887 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7890 = _T_7884 | _T_7889; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7900 = _T_4167 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7901 = _GEN_797 == 7'h7a; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7903 = _T_7901 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7905 = _T_7903 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7906 = _T_7900 | _T_7905; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7916 = _T_4171 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7917 = _GEN_797 == 7'h7b; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7919 = _T_7917 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7921 = _T_7919 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7922 = _T_7916 | _T_7921; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7932 = _T_4175 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7933 = _GEN_797 == 7'h7c; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7935 = _T_7933 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7937 = _T_7935 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7938 = _T_7932 | _T_7937; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7948 = _T_4179 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7949 = _GEN_797 == 7'h7d; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7951 = _T_7949 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7953 = _T_7951 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7954 = _T_7948 | _T_7953; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7964 = _T_4183 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7965 = _GEN_797 == 7'h7e; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7967 = _T_7965 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7969 = _T_7967 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7970 = _T_7964 | _T_7969; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7980 = _T_4187 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7981 = _GEN_797 == 7'h7f; // @[el2_ifu_mem_ctl.scala 754:101]
  wire  _T_7983 = _T_7981 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_7985 = _T_7983 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_7986 = _T_7980 | _T_7985; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_7996 = _T_4063 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_7999 = _T_7485 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8001 = _T_7999 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8002 = _T_7996 | _T_8001; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8012 = _T_4067 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8015 = _T_7501 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8017 = _T_8015 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8018 = _T_8012 | _T_8017; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8028 = _T_4071 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8031 = _T_7517 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8033 = _T_8031 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8034 = _T_8028 | _T_8033; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8044 = _T_4075 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8047 = _T_7533 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8049 = _T_8047 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8050 = _T_8044 | _T_8049; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8060 = _T_4079 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8063 = _T_7549 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8065 = _T_8063 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8066 = _T_8060 | _T_8065; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8076 = _T_4083 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8079 = _T_7565 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8081 = _T_8079 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8082 = _T_8076 | _T_8081; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8092 = _T_4087 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8095 = _T_7581 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8097 = _T_8095 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8098 = _T_8092 | _T_8097; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8108 = _T_4091 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8111 = _T_7597 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8113 = _T_8111 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8114 = _T_8108 | _T_8113; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8124 = _T_4095 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8127 = _T_7613 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8129 = _T_8127 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8130 = _T_8124 | _T_8129; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8140 = _T_4099 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8143 = _T_7629 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8145 = _T_8143 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8146 = _T_8140 | _T_8145; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8156 = _T_4103 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8159 = _T_7645 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8161 = _T_8159 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8162 = _T_8156 | _T_8161; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8172 = _T_4107 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8175 = _T_7661 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8177 = _T_8175 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8178 = _T_8172 | _T_8177; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8188 = _T_4111 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8191 = _T_7677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8193 = _T_8191 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8194 = _T_8188 | _T_8193; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8204 = _T_4115 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8207 = _T_7693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8209 = _T_8207 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8210 = _T_8204 | _T_8209; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8220 = _T_4119 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8223 = _T_7709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8225 = _T_8223 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8226 = _T_8220 | _T_8225; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8236 = _T_4123 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8239 = _T_7725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8241 = _T_8239 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8242 = _T_8236 | _T_8241; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8252 = _T_4127 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8255 = _T_7741 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8257 = _T_8255 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8258 = _T_8252 | _T_8257; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8268 = _T_4131 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8271 = _T_7757 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8273 = _T_8271 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8274 = _T_8268 | _T_8273; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8284 = _T_4135 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8287 = _T_7773 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8289 = _T_8287 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8290 = _T_8284 | _T_8289; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8300 = _T_4139 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8303 = _T_7789 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8305 = _T_8303 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8306 = _T_8300 | _T_8305; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8316 = _T_4143 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8319 = _T_7805 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8321 = _T_8319 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8322 = _T_8316 | _T_8321; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8332 = _T_4147 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8335 = _T_7821 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8337 = _T_8335 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8338 = _T_8332 | _T_8337; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8348 = _T_4151 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8351 = _T_7837 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8353 = _T_8351 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8354 = _T_8348 | _T_8353; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8364 = _T_4155 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8367 = _T_7853 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8369 = _T_8367 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8370 = _T_8364 | _T_8369; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8380 = _T_4159 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8383 = _T_7869 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8385 = _T_8383 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8386 = _T_8380 | _T_8385; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8396 = _T_4163 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8399 = _T_7885 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8401 = _T_8399 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8402 = _T_8396 | _T_8401; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8412 = _T_4167 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8415 = _T_7901 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8417 = _T_8415 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8418 = _T_8412 | _T_8417; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8428 = _T_4171 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8431 = _T_7917 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8433 = _T_8431 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8434 = _T_8428 | _T_8433; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8444 = _T_4175 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8447 = _T_7933 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8449 = _T_8447 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8450 = _T_8444 | _T_8449; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8460 = _T_4179 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8463 = _T_7949 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8465 = _T_8463 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8466 = _T_8460 | _T_8465; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8476 = _T_4183 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8479 = _T_7965 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8481 = _T_8479 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8482 = _T_8476 | _T_8481; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_8492 = _T_4187 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:58]
  wire  _T_8495 = _T_7981 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 754:123]
  wire  _T_8497 = _T_8495 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 754:144]
  wire  _T_8498 = _T_8492 | _T_8497; // @[el2_ifu_mem_ctl.scala 754:80]
  wire  _T_9299 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 808:63]
  wire  _T_9300 = _T_9299 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 808:85]
  wire [1:0] _T_9302 = _T_9300 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9309; // @[el2_ifu_mem_ctl.scala 813:57]
  reg  _T_9310; // @[el2_ifu_mem_ctl.scala 814:56]
  reg  _T_9311; // @[el2_ifu_mem_ctl.scala 815:59]
  wire  _T_9312 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 816:80]
  wire  _T_9313 = ifu_bus_arvalid_ff & _T_9312; // @[el2_ifu_mem_ctl.scala 816:78]
  wire  _T_9314 = _T_9313 & miss_pending; // @[el2_ifu_mem_ctl.scala 816:100]
  reg  _T_9315; // @[el2_ifu_mem_ctl.scala 816:58]
  reg  _T_9316; // @[el2_ifu_mem_ctl.scala 817:58]
  wire  _T_9319 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 824:71]
  wire  _T_9321 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 824:124]
  wire  _T_9323 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 825:50]
  wire  _T_9325 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 825:103]
  wire [3:0] _T_9328 = {_T_9319,_T_9321,_T_9323,_T_9325}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 827:53]
  reg  _T_9339; // @[Reg.scala 27:20]
  rvecc_encode_64 m1 ( // @[el2_ifu_mem_ctl.scala 342:18]
    .io_din(m1_io_din),
    .io_ecc_out(m1_io_ecc_out)
  );
  rvecc_encode_64 m2 ( // @[el2_ifu_mem_ctl.scala 343:18]
    .io_din(m2_io_din),
    .io_ecc_out(m2_io_ecc_out)
  );
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 328:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 327:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 191:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3134; // @[el2_ifu_mem_ctl.scala 704:21]
  assign io_ifu_pmu_ic_miss = _T_9309; // @[el2_ifu_mem_ctl.scala 813:22]
  assign io_ifu_pmu_ic_hit = _T_9310; // @[el2_ifu_mem_ctl.scala 814:21]
  assign io_ifu_pmu_bus_error = _T_9311; // @[el2_ifu_mem_ctl.scala 815:24]
  assign io_ifu_pmu_bus_busy = _T_9315; // @[el2_ifu_mem_ctl.scala 816:23]
  assign io_ifu_pmu_bus_trxn = _T_9316; // @[el2_ifu_mem_ctl.scala 817:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 141:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 140:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 135:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 139:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 137:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 148:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 150:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 145:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 143:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 136:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 134:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 132:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 133:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 142:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 151:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 146:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 566:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_1728; // @[el2_ifu_mem_ctl.scala 567:19]
  assign io_ifu_axi_araddr = _T_1730 & _T_1732; // @[el2_ifu_mem_ctl.scala 568:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 571:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 147:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 569:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 572:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 138:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 570:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 149:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 144:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 573:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 663:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 661:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 665:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 656:20]
  assign io_iccm_ready = _T_1831 & _T_1825; // @[el2_ifu_mem_ctl.scala 636:17]
  assign io_ic_rw_addr = _T_338 | _T_339; // @[el2_ifu_mem_ctl.scala 337:17]
  assign io_ic_wr_en = 2'h0; // @[el2_ifu_mem_ctl.scala 703:15]
  assign io_ic_rd_en = _T_3112 | _T_3117; // @[el2_ifu_mem_ctl.scala 694:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 350:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 350:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 351:23]
  assign io_ifu_ic_debug_rd_data = _T_365; // @[el2_ifu_mem_ctl.scala 359:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 820:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 822:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 823:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 821:25]
  assign io_ic_debug_way = _T_9328[1:0]; // @[el2_ifu_mem_ctl.scala 824:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9302; // @[el2_ifu_mem_ctl.scala 808:19]
  assign io_iccm_rw_addr = _T_2266[14:0]; // @[el2_ifu_mem_ctl.scala 667:19]
  assign io_iccm_wren = _T_1835 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 638:16]
  assign io_iccm_rden = _T_1839 | _T_1840; // @[el2_ifu_mem_ctl.scala 639:16]
  assign io_iccm_wr_data = _T_2241 ? _T_2242 : _T_2249; // @[el2_ifu_mem_ctl.scala 644:19]
  assign io_iccm_wr_size = _T_1845 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 641:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 289:15]
  assign io_ic_access_fault_f = _T_1613 & _T_317; // @[el2_ifu_mem_ctl.scala 391:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_427; // @[el2_ifu_mem_ctl.scala 392:29]
  assign io_iccm_rd_ecc_single_err = _T_3057 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 680:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 681:29]
  assign io_ic_error_start = _T_353 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 353:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 190:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 189:24]
  assign io_ic_fetch_val_f = {_T_435,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 395:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 388:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 385:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 386:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_9339; // @[el2_ifu_mem_ctl.scala 831:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_1618; // @[el2_ifu_mem_ctl.scala 485:27]
  assign io_iccm_correction_state = _T_1646 ? 1'h0 : _GEN_60; // @[el2_ifu_mem_ctl.scala 520:28 el2_ifu_mem_ctl.scala 533:32 el2_ifu_mem_ctl.scala 540:32 el2_ifu_mem_ctl.scala 547:32]
  assign m1_io_din = ifu_bus_rdata_ff; // @[el2_ifu_mem_ctl.scala 344:13]
  assign m2_io_din = {_T_1529,_T_1609}; // @[el2_ifu_mem_ctl.scala 347:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_4322 = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  _T_3678 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_3674 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_3670 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_3666 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_3662 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_3658 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_3654 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_3650 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_3646 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_3642 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_3638 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_3634 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_3630 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_3626 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_3622 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_3618 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_3614 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_3610 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_3606 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_3602 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_3598 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_3594 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_3590 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_3586 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_3582 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_3578 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_3574 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_3570 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_3566 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_3562 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_3558 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_3554 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_3550 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_3546 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_3542 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_3538 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_3534 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_3530 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_3526 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_3522 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_3518 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_3514 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_3510 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_3506 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_3502 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_3498 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_3494 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_3490 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_3486 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_3482 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_3478 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_3474 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_3470 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_3466 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_3462 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_3458 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_3454 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_3450 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_3446 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_3442 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_3438 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_3434 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_3430 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_3426 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_3422 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_3418 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_3414 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_3410 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_3406 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_3402 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_3398 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_3394 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_3390 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_3386 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_3382 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_3378 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_3374 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_3370 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_3366 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_3362 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_3358 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_3354 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_3350 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_3346 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_3342 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_3338 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_3334 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_3330 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_3326 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_3322 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_3318 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_3314 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_3310 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_3306 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_3302 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_3298 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_3294 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_3290 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_3286 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_3282 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_3278 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_3274 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_3270 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_3266 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_3262 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_3258 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_3254 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_3250 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_3246 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_3242 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_3238 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_3234 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_3230 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_3226 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_3222 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_3218 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_3214 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_3210 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3206 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3202 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3198 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3194 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3190 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3186 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3182 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3178 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  _T_3174 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _T_3170 = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_151[30:0];
  _RAND_152 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  reset_ic_ff = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  miss_addr = _RAND_159[25:0];
  _RAND_160 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_161[2:0];
  _RAND_162 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_162[0:0];
  _RAND_163 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_163[63:0];
  _RAND_164 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_440[0:0];
  _RAND_441 = {3{`RANDOM}};
  _T_365 = _RAND_441[70:0];
  _RAND_442 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_445[2:0];
  _RAND_446 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_448[0:0];
  _RAND_449 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_449[38:0];
  _RAND_450 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_451[2:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_453[0:0];
  _RAND_454 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_454[63:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_455[13:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_457[13:0];
  _RAND_458 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_458[6:0];
  _RAND_459 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_new_ff = _RAND_460[2:0];
  _RAND_461 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  ic_valid_ff = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_9309 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_9310 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_9311 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_9315 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_9316 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_9339 = _RAND_468[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      _T_3678 <= 3'h0;
    end else if (_T_3677) begin
      _T_3678 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3674 <= 3'h0;
    end else if (_T_3673) begin
      _T_3674 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3670 <= 3'h0;
    end else if (_T_3669) begin
      _T_3670 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3666 <= 3'h0;
    end else if (_T_3665) begin
      _T_3666 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3662 <= 3'h0;
    end else if (_T_3661) begin
      _T_3662 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3658 <= 3'h0;
    end else if (_T_3657) begin
      _T_3658 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3654 <= 3'h0;
    end else if (_T_3653) begin
      _T_3654 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3650 <= 3'h0;
    end else if (_T_3649) begin
      _T_3650 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3646 <= 3'h0;
    end else if (_T_3645) begin
      _T_3646 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3642 <= 3'h0;
    end else if (_T_3641) begin
      _T_3642 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3638 <= 3'h0;
    end else if (_T_3637) begin
      _T_3638 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3634 <= 3'h0;
    end else if (_T_3633) begin
      _T_3634 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3630 <= 3'h0;
    end else if (_T_3629) begin
      _T_3630 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3626 <= 3'h0;
    end else if (_T_3625) begin
      _T_3626 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3622 <= 3'h0;
    end else if (_T_3621) begin
      _T_3622 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3618 <= 3'h0;
    end else if (_T_3617) begin
      _T_3618 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3614 <= 3'h0;
    end else if (_T_3613) begin
      _T_3614 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3610 <= 3'h0;
    end else if (_T_3609) begin
      _T_3610 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3606 <= 3'h0;
    end else if (_T_3605) begin
      _T_3606 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3602 <= 3'h0;
    end else if (_T_3601) begin
      _T_3602 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3598 <= 3'h0;
    end else if (_T_3597) begin
      _T_3598 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3594 <= 3'h0;
    end else if (_T_3593) begin
      _T_3594 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3590 <= 3'h0;
    end else if (_T_3589) begin
      _T_3590 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3586 <= 3'h0;
    end else if (_T_3585) begin
      _T_3586 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3582 <= 3'h0;
    end else if (_T_3581) begin
      _T_3582 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3578 <= 3'h0;
    end else if (_T_3577) begin
      _T_3578 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3574 <= 3'h0;
    end else if (_T_3573) begin
      _T_3574 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3570 <= 3'h0;
    end else if (_T_3569) begin
      _T_3570 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3566 <= 3'h0;
    end else if (_T_3565) begin
      _T_3566 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3562 <= 3'h0;
    end else if (_T_3561) begin
      _T_3562 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3558 <= 3'h0;
    end else if (_T_3557) begin
      _T_3558 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3554 <= 3'h0;
    end else if (_T_3553) begin
      _T_3554 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3550 <= 3'h0;
    end else if (_T_3549) begin
      _T_3550 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3546 <= 3'h0;
    end else if (_T_3545) begin
      _T_3546 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3542 <= 3'h0;
    end else if (_T_3541) begin
      _T_3542 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3538 <= 3'h0;
    end else if (_T_3537) begin
      _T_3538 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3534 <= 3'h0;
    end else if (_T_3533) begin
      _T_3534 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3530 <= 3'h0;
    end else if (_T_3529) begin
      _T_3530 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3526 <= 3'h0;
    end else if (_T_3525) begin
      _T_3526 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3522 <= 3'h0;
    end else if (_T_3521) begin
      _T_3522 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3518 <= 3'h0;
    end else if (_T_3517) begin
      _T_3518 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3514 <= 3'h0;
    end else if (_T_3513) begin
      _T_3514 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3510 <= 3'h0;
    end else if (_T_3509) begin
      _T_3510 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3506 <= 3'h0;
    end else if (_T_3505) begin
      _T_3506 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3502 <= 3'h0;
    end else if (_T_3501) begin
      _T_3502 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3498 <= 3'h0;
    end else if (_T_3497) begin
      _T_3498 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3494 <= 3'h0;
    end else if (_T_3493) begin
      _T_3494 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3490 <= 3'h0;
    end else if (_T_3489) begin
      _T_3490 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3486 <= 3'h0;
    end else if (_T_3485) begin
      _T_3486 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3482 <= 3'h0;
    end else if (_T_3481) begin
      _T_3482 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3478 <= 3'h0;
    end else if (_T_3477) begin
      _T_3478 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3474 <= 3'h0;
    end else if (_T_3473) begin
      _T_3474 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3470 <= 3'h0;
    end else if (_T_3469) begin
      _T_3470 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3466 <= 3'h0;
    end else if (_T_3465) begin
      _T_3466 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3462 <= 3'h0;
    end else if (_T_3461) begin
      _T_3462 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3458 <= 3'h0;
    end else if (_T_3457) begin
      _T_3458 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3454 <= 3'h0;
    end else if (_T_3453) begin
      _T_3454 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3450 <= 3'h0;
    end else if (_T_3449) begin
      _T_3450 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3446 <= 3'h0;
    end else if (_T_3445) begin
      _T_3446 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3442 <= 3'h0;
    end else if (_T_3441) begin
      _T_3442 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3438 <= 3'h0;
    end else if (_T_3437) begin
      _T_3438 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3434 <= 3'h0;
    end else if (_T_3433) begin
      _T_3434 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3430 <= 3'h0;
    end else if (_T_3429) begin
      _T_3430 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3426 <= 3'h0;
    end else if (_T_3425) begin
      _T_3426 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3422 <= 3'h0;
    end else if (_T_3421) begin
      _T_3422 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3418 <= 3'h0;
    end else if (_T_3417) begin
      _T_3418 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3414 <= 3'h0;
    end else if (_T_3413) begin
      _T_3414 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3410 <= 3'h0;
    end else if (_T_3409) begin
      _T_3410 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3406 <= 3'h0;
    end else if (_T_3405) begin
      _T_3406 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3402 <= 3'h0;
    end else if (_T_3401) begin
      _T_3402 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3398 <= 3'h0;
    end else if (_T_3397) begin
      _T_3398 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3394 <= 3'h0;
    end else if (_T_3393) begin
      _T_3394 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3390 <= 3'h0;
    end else if (_T_3389) begin
      _T_3390 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3386 <= 3'h0;
    end else if (_T_3385) begin
      _T_3386 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3382 <= 3'h0;
    end else if (_T_3381) begin
      _T_3382 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3378 <= 3'h0;
    end else if (_T_3377) begin
      _T_3378 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3374 <= 3'h0;
    end else if (_T_3373) begin
      _T_3374 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3370 <= 3'h0;
    end else if (_T_3369) begin
      _T_3370 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3366 <= 3'h0;
    end else if (_T_3365) begin
      _T_3366 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3362 <= 3'h0;
    end else if (_T_3361) begin
      _T_3362 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3358 <= 3'h0;
    end else if (_T_3357) begin
      _T_3358 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3354 <= 3'h0;
    end else if (_T_3353) begin
      _T_3354 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3350 <= 3'h0;
    end else if (_T_3349) begin
      _T_3350 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3346 <= 3'h0;
    end else if (_T_3345) begin
      _T_3346 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3342 <= 3'h0;
    end else if (_T_3341) begin
      _T_3342 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3338 <= 3'h0;
    end else if (_T_3337) begin
      _T_3338 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3334 <= 3'h0;
    end else if (_T_3333) begin
      _T_3334 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3330 <= 3'h0;
    end else if (_T_3329) begin
      _T_3330 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3326 <= 3'h0;
    end else if (_T_3325) begin
      _T_3326 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3322 <= 3'h0;
    end else if (_T_3321) begin
      _T_3322 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3318 <= 3'h0;
    end else if (_T_3317) begin
      _T_3318 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3314 <= 3'h0;
    end else if (_T_3313) begin
      _T_3314 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3310 <= 3'h0;
    end else if (_T_3309) begin
      _T_3310 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3306 <= 3'h0;
    end else if (_T_3305) begin
      _T_3306 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3302 <= 3'h0;
    end else if (_T_3301) begin
      _T_3302 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3298 <= 3'h0;
    end else if (_T_3297) begin
      _T_3298 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3294 <= 3'h0;
    end else if (_T_3293) begin
      _T_3294 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3290 <= 3'h0;
    end else if (_T_3289) begin
      _T_3290 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3286 <= 3'h0;
    end else if (_T_3285) begin
      _T_3286 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3282 <= 3'h0;
    end else if (_T_3281) begin
      _T_3282 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3278 <= 3'h0;
    end else if (_T_3277) begin
      _T_3278 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3274 <= 3'h0;
    end else if (_T_3273) begin
      _T_3274 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3270 <= 3'h0;
    end else if (_T_3269) begin
      _T_3270 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3266 <= 3'h0;
    end else if (_T_3265) begin
      _T_3266 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3262 <= 3'h0;
    end else if (_T_3261) begin
      _T_3262 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3258 <= 3'h0;
    end else if (_T_3257) begin
      _T_3258 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3254 <= 3'h0;
    end else if (_T_3253) begin
      _T_3254 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3250 <= 3'h0;
    end else if (_T_3249) begin
      _T_3250 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3246 <= 3'h0;
    end else if (_T_3245) begin
      _T_3246 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3242 <= 3'h0;
    end else if (_T_3241) begin
      _T_3242 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3238 <= 3'h0;
    end else if (_T_3237) begin
      _T_3238 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3234 <= 3'h0;
    end else if (_T_3233) begin
      _T_3234 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3230 <= 3'h0;
    end else if (_T_3229) begin
      _T_3230 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3226 <= 3'h0;
    end else if (_T_3225) begin
      _T_3226 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3222 <= 3'h0;
    end else if (_T_3221) begin
      _T_3222 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3218 <= 3'h0;
    end else if (_T_3217) begin
      _T_3218 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3214 <= 3'h0;
    end else if (_T_3213) begin
      _T_3214 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3210 <= 3'h0;
    end else if (_T_3209) begin
      _T_3210 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3206 <= 3'h0;
    end else if (_T_3205) begin
      _T_3206 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3202 <= 3'h0;
    end else if (_T_3201) begin
      _T_3202 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3198 <= 3'h0;
    end else if (_T_3197) begin
      _T_3198 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3194 <= 3'h0;
    end else if (_T_3193) begin
      _T_3194 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3190 <= 3'h0;
    end else if (_T_3189) begin
      _T_3190 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3186 <= 3'h0;
    end else if (_T_3185) begin
      _T_3186 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3182 <= 3'h0;
    end else if (_T_3181) begin
      _T_3182 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3178 <= 3'h0;
    end else if (_T_3177) begin
      _T_3178 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3174 <= 3'h0;
    end else if (_T_3173) begin
      _T_3174 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3170 <= 3'h0;
    end else if (_T_3169) begin
      _T_3170 <= way_status_new_ff;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_289;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= 2'h0;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_1771) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_1767;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_4930) begin
      ic_tag_valid_out_1_0 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_4946) begin
      ic_tag_valid_out_1_1 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_4962) begin
      ic_tag_valid_out_1_2 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_4978) begin
      ic_tag_valid_out_1_3 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_4994) begin
      ic_tag_valid_out_1_4 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5010) begin
      ic_tag_valid_out_1_5 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5026) begin
      ic_tag_valid_out_1_6 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5042) begin
      ic_tag_valid_out_1_7 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5058) begin
      ic_tag_valid_out_1_8 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5074) begin
      ic_tag_valid_out_1_9 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5090) begin
      ic_tag_valid_out_1_10 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5106) begin
      ic_tag_valid_out_1_11 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5122) begin
      ic_tag_valid_out_1_12 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5138) begin
      ic_tag_valid_out_1_13 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5154) begin
      ic_tag_valid_out_1_14 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5170) begin
      ic_tag_valid_out_1_15 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5186) begin
      ic_tag_valid_out_1_16 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5202) begin
      ic_tag_valid_out_1_17 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5218) begin
      ic_tag_valid_out_1_18 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5234) begin
      ic_tag_valid_out_1_19 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5250) begin
      ic_tag_valid_out_1_20 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5266) begin
      ic_tag_valid_out_1_21 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5282) begin
      ic_tag_valid_out_1_22 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5298) begin
      ic_tag_valid_out_1_23 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_5314) begin
      ic_tag_valid_out_1_24 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_5330) begin
      ic_tag_valid_out_1_25 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_5346) begin
      ic_tag_valid_out_1_26 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_5362) begin
      ic_tag_valid_out_1_27 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_5378) begin
      ic_tag_valid_out_1_28 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_5394) begin
      ic_tag_valid_out_1_29 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_5410) begin
      ic_tag_valid_out_1_30 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_5426) begin
      ic_tag_valid_out_1_31 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_5954) begin
      ic_tag_valid_out_1_32 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_5970) begin
      ic_tag_valid_out_1_33 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_5986) begin
      ic_tag_valid_out_1_34 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6002) begin
      ic_tag_valid_out_1_35 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6018) begin
      ic_tag_valid_out_1_36 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6034) begin
      ic_tag_valid_out_1_37 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6050) begin
      ic_tag_valid_out_1_38 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6066) begin
      ic_tag_valid_out_1_39 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6082) begin
      ic_tag_valid_out_1_40 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6098) begin
      ic_tag_valid_out_1_41 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6114) begin
      ic_tag_valid_out_1_42 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6130) begin
      ic_tag_valid_out_1_43 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6146) begin
      ic_tag_valid_out_1_44 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6162) begin
      ic_tag_valid_out_1_45 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6178) begin
      ic_tag_valid_out_1_46 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6194) begin
      ic_tag_valid_out_1_47 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6210) begin
      ic_tag_valid_out_1_48 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6226) begin
      ic_tag_valid_out_1_49 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6242) begin
      ic_tag_valid_out_1_50 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6258) begin
      ic_tag_valid_out_1_51 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6274) begin
      ic_tag_valid_out_1_52 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6290) begin
      ic_tag_valid_out_1_53 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6306) begin
      ic_tag_valid_out_1_54 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6322) begin
      ic_tag_valid_out_1_55 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6338) begin
      ic_tag_valid_out_1_56 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6354) begin
      ic_tag_valid_out_1_57 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6370) begin
      ic_tag_valid_out_1_58 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_6386) begin
      ic_tag_valid_out_1_59 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_6402) begin
      ic_tag_valid_out_1_60 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_6418) begin
      ic_tag_valid_out_1_61 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_6434) begin
      ic_tag_valid_out_1_62 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_6450) begin
      ic_tag_valid_out_1_63 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_6978) begin
      ic_tag_valid_out_1_64 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_6994) begin
      ic_tag_valid_out_1_65 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7010) begin
      ic_tag_valid_out_1_66 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7026) begin
      ic_tag_valid_out_1_67 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7042) begin
      ic_tag_valid_out_1_68 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7058) begin
      ic_tag_valid_out_1_69 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7074) begin
      ic_tag_valid_out_1_70 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7090) begin
      ic_tag_valid_out_1_71 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7106) begin
      ic_tag_valid_out_1_72 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7122) begin
      ic_tag_valid_out_1_73 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7138) begin
      ic_tag_valid_out_1_74 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7154) begin
      ic_tag_valid_out_1_75 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7170) begin
      ic_tag_valid_out_1_76 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7186) begin
      ic_tag_valid_out_1_77 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7202) begin
      ic_tag_valid_out_1_78 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7218) begin
      ic_tag_valid_out_1_79 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7234) begin
      ic_tag_valid_out_1_80 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7250) begin
      ic_tag_valid_out_1_81 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7266) begin
      ic_tag_valid_out_1_82 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7282) begin
      ic_tag_valid_out_1_83 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7298) begin
      ic_tag_valid_out_1_84 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7314) begin
      ic_tag_valid_out_1_85 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7330) begin
      ic_tag_valid_out_1_86 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7346) begin
      ic_tag_valid_out_1_87 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7362) begin
      ic_tag_valid_out_1_88 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7378) begin
      ic_tag_valid_out_1_89 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7394) begin
      ic_tag_valid_out_1_90 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7410) begin
      ic_tag_valid_out_1_91 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7426) begin
      ic_tag_valid_out_1_92 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7442) begin
      ic_tag_valid_out_1_93 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_7458) begin
      ic_tag_valid_out_1_94 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_7474) begin
      ic_tag_valid_out_1_95 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8002) begin
      ic_tag_valid_out_1_96 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8018) begin
      ic_tag_valid_out_1_97 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8034) begin
      ic_tag_valid_out_1_98 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8050) begin
      ic_tag_valid_out_1_99 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8066) begin
      ic_tag_valid_out_1_100 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8082) begin
      ic_tag_valid_out_1_101 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8098) begin
      ic_tag_valid_out_1_102 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8114) begin
      ic_tag_valid_out_1_103 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8130) begin
      ic_tag_valid_out_1_104 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8146) begin
      ic_tag_valid_out_1_105 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8162) begin
      ic_tag_valid_out_1_106 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8178) begin
      ic_tag_valid_out_1_107 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8194) begin
      ic_tag_valid_out_1_108 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8210) begin
      ic_tag_valid_out_1_109 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8226) begin
      ic_tag_valid_out_1_110 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8242) begin
      ic_tag_valid_out_1_111 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8258) begin
      ic_tag_valid_out_1_112 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8274) begin
      ic_tag_valid_out_1_113 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8290) begin
      ic_tag_valid_out_1_114 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8306) begin
      ic_tag_valid_out_1_115 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8322) begin
      ic_tag_valid_out_1_116 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8338) begin
      ic_tag_valid_out_1_117 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8354) begin
      ic_tag_valid_out_1_118 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8370) begin
      ic_tag_valid_out_1_119 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8386) begin
      ic_tag_valid_out_1_120 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8402) begin
      ic_tag_valid_out_1_121 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8418) begin
      ic_tag_valid_out_1_122 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8434) begin
      ic_tag_valid_out_1_123 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8450) begin
      ic_tag_valid_out_1_124 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8466) begin
      ic_tag_valid_out_1_125 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8482) begin
      ic_tag_valid_out_1_126 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8498) begin
      ic_tag_valid_out_1_127 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_4418) begin
      ic_tag_valid_out_0_0 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_4434) begin
      ic_tag_valid_out_0_1 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_4450) begin
      ic_tag_valid_out_0_2 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_4466) begin
      ic_tag_valid_out_0_3 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_4482) begin
      ic_tag_valid_out_0_4 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_4498) begin
      ic_tag_valid_out_0_5 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_4514) begin
      ic_tag_valid_out_0_6 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_4530) begin
      ic_tag_valid_out_0_7 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_4546) begin
      ic_tag_valid_out_0_8 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_4562) begin
      ic_tag_valid_out_0_9 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_4578) begin
      ic_tag_valid_out_0_10 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_4594) begin
      ic_tag_valid_out_0_11 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_4610) begin
      ic_tag_valid_out_0_12 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_4626) begin
      ic_tag_valid_out_0_13 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_4642) begin
      ic_tag_valid_out_0_14 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_4658) begin
      ic_tag_valid_out_0_15 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_4674) begin
      ic_tag_valid_out_0_16 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_4690) begin
      ic_tag_valid_out_0_17 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_4706) begin
      ic_tag_valid_out_0_18 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_4722) begin
      ic_tag_valid_out_0_19 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_4738) begin
      ic_tag_valid_out_0_20 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_4754) begin
      ic_tag_valid_out_0_21 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_4770) begin
      ic_tag_valid_out_0_22 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_4786) begin
      ic_tag_valid_out_0_23 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_4802) begin
      ic_tag_valid_out_0_24 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_4818) begin
      ic_tag_valid_out_0_25 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_4834) begin
      ic_tag_valid_out_0_26 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_4850) begin
      ic_tag_valid_out_0_27 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_4866) begin
      ic_tag_valid_out_0_28 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_4882) begin
      ic_tag_valid_out_0_29 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_4898) begin
      ic_tag_valid_out_0_30 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_4914) begin
      ic_tag_valid_out_0_31 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_5442) begin
      ic_tag_valid_out_0_32 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_5458) begin
      ic_tag_valid_out_0_33 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_5474) begin
      ic_tag_valid_out_0_34 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_5490) begin
      ic_tag_valid_out_0_35 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_5506) begin
      ic_tag_valid_out_0_36 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_5522) begin
      ic_tag_valid_out_0_37 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_5538) begin
      ic_tag_valid_out_0_38 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_5554) begin
      ic_tag_valid_out_0_39 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_5570) begin
      ic_tag_valid_out_0_40 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_5586) begin
      ic_tag_valid_out_0_41 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_5602) begin
      ic_tag_valid_out_0_42 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_5618) begin
      ic_tag_valid_out_0_43 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_5634) begin
      ic_tag_valid_out_0_44 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_5650) begin
      ic_tag_valid_out_0_45 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_5666) begin
      ic_tag_valid_out_0_46 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_5682) begin
      ic_tag_valid_out_0_47 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_5698) begin
      ic_tag_valid_out_0_48 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_5714) begin
      ic_tag_valid_out_0_49 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_5730) begin
      ic_tag_valid_out_0_50 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_5746) begin
      ic_tag_valid_out_0_51 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_5762) begin
      ic_tag_valid_out_0_52 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_5778) begin
      ic_tag_valid_out_0_53 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_5794) begin
      ic_tag_valid_out_0_54 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_5810) begin
      ic_tag_valid_out_0_55 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_5826) begin
      ic_tag_valid_out_0_56 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_5842) begin
      ic_tag_valid_out_0_57 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_5858) begin
      ic_tag_valid_out_0_58 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_5874) begin
      ic_tag_valid_out_0_59 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_5890) begin
      ic_tag_valid_out_0_60 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_5906) begin
      ic_tag_valid_out_0_61 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_5922) begin
      ic_tag_valid_out_0_62 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_5938) begin
      ic_tag_valid_out_0_63 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_6466) begin
      ic_tag_valid_out_0_64 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_6482) begin
      ic_tag_valid_out_0_65 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_6498) begin
      ic_tag_valid_out_0_66 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_6514) begin
      ic_tag_valid_out_0_67 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_6530) begin
      ic_tag_valid_out_0_68 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_6546) begin
      ic_tag_valid_out_0_69 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_6562) begin
      ic_tag_valid_out_0_70 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_6578) begin
      ic_tag_valid_out_0_71 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_6594) begin
      ic_tag_valid_out_0_72 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_6610) begin
      ic_tag_valid_out_0_73 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_6626) begin
      ic_tag_valid_out_0_74 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_6642) begin
      ic_tag_valid_out_0_75 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_6658) begin
      ic_tag_valid_out_0_76 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_6674) begin
      ic_tag_valid_out_0_77 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_6690) begin
      ic_tag_valid_out_0_78 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_6706) begin
      ic_tag_valid_out_0_79 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_6722) begin
      ic_tag_valid_out_0_80 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_6738) begin
      ic_tag_valid_out_0_81 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_6754) begin
      ic_tag_valid_out_0_82 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_6770) begin
      ic_tag_valid_out_0_83 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_6786) begin
      ic_tag_valid_out_0_84 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_6802) begin
      ic_tag_valid_out_0_85 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_6818) begin
      ic_tag_valid_out_0_86 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_6834) begin
      ic_tag_valid_out_0_87 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_6850) begin
      ic_tag_valid_out_0_88 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_6866) begin
      ic_tag_valid_out_0_89 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_6882) begin
      ic_tag_valid_out_0_90 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_6898) begin
      ic_tag_valid_out_0_91 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_6914) begin
      ic_tag_valid_out_0_92 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_6930) begin
      ic_tag_valid_out_0_93 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_6946) begin
      ic_tag_valid_out_0_94 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_6962) begin
      ic_tag_valid_out_0_95 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_7490) begin
      ic_tag_valid_out_0_96 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_7506) begin
      ic_tag_valid_out_0_97 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_7522) begin
      ic_tag_valid_out_0_98 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_7538) begin
      ic_tag_valid_out_0_99 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_7554) begin
      ic_tag_valid_out_0_100 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_7570) begin
      ic_tag_valid_out_0_101 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_7586) begin
      ic_tag_valid_out_0_102 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_7602) begin
      ic_tag_valid_out_0_103 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_7618) begin
      ic_tag_valid_out_0_104 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_7634) begin
      ic_tag_valid_out_0_105 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_7650) begin
      ic_tag_valid_out_0_106 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_7666) begin
      ic_tag_valid_out_0_107 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_7682) begin
      ic_tag_valid_out_0_108 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_7698) begin
      ic_tag_valid_out_0_109 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_7714) begin
      ic_tag_valid_out_0_110 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_7730) begin
      ic_tag_valid_out_0_111 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_7746) begin
      ic_tag_valid_out_0_112 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_7762) begin
      ic_tag_valid_out_0_113 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_7778) begin
      ic_tag_valid_out_0_114 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_7794) begin
      ic_tag_valid_out_0_115 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_7810) begin
      ic_tag_valid_out_0_116 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_7826) begin
      ic_tag_valid_out_0_117 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_7842) begin
      ic_tag_valid_out_0_118 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_7858) begin
      ic_tag_valid_out_0_119 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_7874) begin
      ic_tag_valid_out_0_120 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_7890) begin
      ic_tag_valid_out_0_121 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_7906) begin
      ic_tag_valid_out_0_122 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_7922) begin
      ic_tag_valid_out_0_123 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_7938) begin
      ic_tag_valid_out_0_124 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_7954) begin
      ic_tag_valid_out_0_125 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_7970) begin
      ic_tag_valid_out_0_126 <= _T_4409;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_7986) begin
      ic_tag_valid_out_0_127 <= _T_4409;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_365 <= 71'h0;
    end else if (ic_debug_rd_en_ff) begin
      if (ic_debug_ict_array_sel_ff) begin
        _T_365 <= {{5'd0}, _T_364};
      end else begin
        _T_365 <= io_ic_debug_rd_data;
      end
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_1720) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_1795) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_1839;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_1621) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_1623) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_1633) begin
        perr_state <= 3'h0;
      end else if (_T_1636) begin
        if (_T_1638) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_1642) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_1646) begin
        err_stop_state <= 2'h1;
      end else if (_T_1651) begin
        if (_T_1653) begin
          err_stop_state <= 2'h0;
        end else if (_T_1674) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_1678) begin
        if (_T_1653) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_1695) begin
        if (_T_1699) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_524;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_4322 <= 7'h0;
    end else if (_T_3143) begin
      _T_4322 <= io_ic_debug_addr[9:3];
    end else begin
      _T_4322 <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_564;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3078;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_2253;
    end else begin
      iccm_dma_rdata <= _T_2254;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3074;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3143) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3146) begin
      way_status_new_ff <= _T_3150;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3146) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_9339 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_9339 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_9309 <= 1'h0;
    end else begin
      _T_9309 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_9310 <= 1'h0;
    end else begin
      _T_9310 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_9311 <= 1'h0;
    end else begin
      _T_9311 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_9315 <= 1'h0;
    end else begin
      _T_9315 <= _T_9314;
    end
    if (reset) begin
      _T_9316 <= 1'h0;
    end else begin
      _T_9316 <= bus_cmd_sent;
    end
  end
endmodule
